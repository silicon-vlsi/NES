magic
tech sky130A
timestamp 1766556303
<< locali >>
rect 181 1714 7509 1722
rect 181 1650 191 1714
rect 359 1650 7509 1714
rect 181 1642 7509 1650
rect -708 1592 1428 1593
rect -708 1512 1944 1592
rect -192 1511 1944 1512
rect -469 1423 -336 1433
rect -469 1352 -457 1423
rect -356 1352 -336 1423
rect -469 -2662 -336 1352
rect 3255 386 3333 460
rect 3269 -441 3381 -361
rect 681 -465 1611 -464
rect 681 -477 1908 -465
rect 70 -483 1908 -477
rect 58 -612 1908 -483
rect 283 -670 1908 -612
rect 3269 -540 3280 -441
rect 3371 -540 3381 -441
rect 283 -679 1611 -670
rect 681 -691 1611 -679
rect 3088 -1336 3208 -1239
rect 3168 -1337 3208 -1336
rect 3269 -1841 3381 -540
rect 8398 -894 8499 -841
rect 3269 -1933 3282 -1841
rect 3369 -1933 3381 -1841
rect 3269 -1945 3381 -1933
rect 3081 -2252 3625 -2035
rect 3080 -2653 3639 -2434
rect -469 -2765 -451 -2662
rect -353 -2765 -336 -2662
rect -469 -2780 -336 -2765
rect 1396 -3017 1687 -2943
<< viali >>
rect 191 1650 359 1714
rect -457 1352 -356 1423
rect 2807 384 2924 461
rect -293 -687 283 -612
rect 3280 -540 3371 -441
rect 3282 -1933 3369 -1841
rect -451 -2765 -353 -2662
<< metal1 >>
rect -468 1722 -335 1723
rect -468 1714 369 1722
rect -468 1650 191 1714
rect 359 1650 369 1714
rect -468 1642 369 1650
rect -468 1423 -335 1642
rect -468 1352 -457 1423
rect -356 1352 -335 1423
rect -468 1345 -335 1352
rect 2798 470 2938 473
rect 2798 461 2939 470
rect 2798 384 2807 461
rect 2924 384 2939 461
rect 1989 -42 2209 -39
rect 1989 -137 2210 -42
rect 1989 -364 2088 -137
rect 2798 -191 2939 384
rect 8561 369 9553 473
rect 9366 332 9618 333
rect 9213 232 9618 332
rect 9271 231 9618 232
rect 2798 -342 3223 -191
rect 9271 -255 9469 231
rect -671 -612 314 -604
rect -671 -687 -293 -612
rect 283 -687 314 -612
rect -671 -696 314 -687
rect 3054 -864 3222 -342
rect 8633 -393 11168 -255
rect 3268 -441 8543 -428
rect 3268 -540 3280 -441
rect 3371 -540 8543 -441
rect 3268 -555 8543 -540
rect 3268 -557 8260 -555
rect 3268 -558 5884 -557
rect 3055 -975 3208 -864
rect 3687 -874 3999 -752
rect 8219 -1574 8320 -1564
rect -677 -1793 195 -1680
rect 3004 -1682 3517 -1681
rect 3004 -1684 3606 -1682
rect 2678 -1696 3606 -1684
rect 2678 -1785 3399 -1696
rect 3540 -1785 3606 -1696
rect 2678 -1796 3606 -1785
rect 3004 -1798 3606 -1796
rect 3004 -1799 3517 -1798
rect -679 -1943 303 -1833
rect 3180 -1841 3379 -1832
rect 3180 -1933 3282 -1841
rect 3369 -1933 3379 -1841
rect 3180 -1943 3379 -1933
rect 3185 -1945 3379 -1943
rect 8219 -1870 8232 -1574
rect 8313 -1870 8320 -1574
rect 8219 -1938 8320 -1870
rect 8219 -2062 8690 -1938
rect 10682 -2060 11450 -1934
rect 8227 -2253 8335 -2239
rect 8227 -2527 8237 -2253
rect 8324 -2527 8335 -2253
rect -467 -2662 -337 -2648
rect -467 -2765 -451 -2662
rect -353 -2765 -337 -2662
rect -467 -2783 -337 -2765
rect -467 -2892 281 -2783
rect -384 -2893 281 -2892
rect 8227 -3275 8335 -2527
rect 8227 -3277 8691 -3275
rect 8227 -3426 11450 -3277
<< via1 >>
rect 3399 -1785 3540 -1696
rect 8232 -1870 8313 -1574
rect 8237 -2527 8324 -2253
<< metal2 >>
rect 3384 -1696 6019 -1573
rect 3384 -1785 3399 -1696
rect 3540 -1785 6019 -1696
rect 3384 -1873 6019 -1785
rect 6375 -1574 8319 -1565
rect 6375 -1870 8232 -1574
rect 8313 -1870 8319 -1574
rect 6375 -1896 8319 -1870
rect 5699 -2241 8337 -2238
rect 5698 -2253 8337 -2241
rect 5698 -2527 8237 -2253
rect 8324 -2527 8337 -2253
rect 5698 -2549 8337 -2527
rect 5698 -2551 8174 -2549
use BGR_bjt_copy  BGR_bjt_copy_0
timestamp 1764841004
transform 1 0 3507 0 1 -2663
box -117 -740 4829 1943
use BGR_nmostrial_copy  BGR_nmostrial_copy_0
timestamp 1766123683
transform 1 0 -18 0 1 -1763
box -300 -1270 3266 1170
use BGR_pmos2  BGR_pmos2_0
timestamp 1766556163
transform 1 0 3809 0 1 792
box -4060 -930 5470 1130
use BGR_resistor_copy  BGR_resistor_copy_0
timestamp 1764841088
transform 1 0 8458 0 1 -1538
box -105 -2050 2597 1450
use BGR_starternmos_copy  BGR_starternmos_copy_0
timestamp 1766122499
transform 1 0 980 0 1 -264
box -930 -270 1040 170
<< labels >>
rlabel space 8064 1550 8064 1550 1 vdd
rlabel locali -655 1547 -655 1547 1 vdd
port 5 n
rlabel metal1 9526 262 9526 262 1 vref
port 10 n
rlabel metal1 -651 -653 -651 -653 1 gnd
port 8 n
<< end >>
