** sch_path: /home/somya/work/xschem/BGR_final_copy_sc.sch
.title BGR-sc  test
*.include /home/somya/sim/BGR_layoutpex.spice
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.temp 27
.global VDD GND

*.PININFO vdd:B vref:B gnd:B gnd:B gnd:B gnd:B gnd:B
XR2 net4 net6 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR1 net4 net6 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR3 net7 net8 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR4 net6 net7 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR5 net9 vref gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR6 net10 net9 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR7 net11 net10 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR8 net21 net11 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR9 net12 net21 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR10 net13 net12 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR11 net14 net13 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR12 net22 net14 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR13 net15 net22 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR14 net16 net15 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR15 net17 net16 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR16 net23 net17 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR17 net18 net23 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR18 net19 net18 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR19 net20 net19 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR20 net24 net20 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR21 net24 net25 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XR22 net24 net25 gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=1 m=1
XRdummy gnd gnd gnd sky130_fd_pr__res_high_po_1p41 L=7.58 mult=4 m=4
XQ4 gnd gnd net8 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=8
XQ5 gnd gnd net25 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
XQ6 gnd gnd net3 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
Xdummy gnd gnd gnd sky130_fd_pr__pnp_05v5_W3p40L3p40 m=18
XM1 net26 net2 vdd VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
XM2 pmosterminal net2 net26 VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
XM4 net1 pmosterminal net2 VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
XM3 net1 net2 vdd VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=4
XM5 net2 net2 vdd VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=4
XM6 vref net2 vdd VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=4
Xpdummy1 net2 vdd vdd VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=5 nf=1 m=1
Xpdummy2 pmosterminal vdd vdd VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=5 nf=1 m=1
Xpdummy3 net2 vdd vdd VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
Xpfldummy4 vdd vdd vdd VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=4
XMN3 net5 net5 gnd GND sky130_fd_pr__nfet_01v8_lvt L=7 W=1 nf=1 m=1
XMN4 pmosterminal pmosterminal net5 GND sky130_fd_pr__nfet_01v8_lvt L=7 W=1 nf=1 m=1
Xndummy1 net4 gnd gnd GND sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 m=4
Xndummy2 net1 gnd gnd GND sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 m=6
Xndummy3 net2 gnd gnd GND sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 m=2
XMN1 net1 net1 net3 GND sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 m=8
XMN2 net2 net1 net4 GND sky130_fd_pr__nfet_01v8_lvt L=1 W=5 nf=1 m=8

*.ends
*** supply voltage
*.dc    vsup    0       3.3     0.3.3

vsup    vdd     gnd     dc      2

.dc temp -40 125 5

*vsup   vdd     gnd     pulse   0       2       10n     1u      1u      1m      100u
*.tran  5n      10u

.control
run
plot v(vref)
*plot vid1#branch vid2#branch vid3#branch vid4#branch vid5#branch

.endc
.end
     
