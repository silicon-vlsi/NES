magic
tech sky130A
timestamp 1766556163
<< nwell >>
rect -4060 930 5150 1130
rect -4060 500 -3830 930
rect 4960 500 5150 930
rect -4060 -200 5150 500
rect -4060 -570 -3830 -200
rect -2150 -300 -1850 -200
rect 4960 -570 5150 -200
rect -4060 -800 5150 -570
<< pmoslvt >>
rect -3550 -100 -3350 400
rect -3150 -100 -2950 400
rect -2700 -100 -2600 400
rect -2400 -100 -2300 400
rect -2100 -100 -2000 400
rect -1850 -100 -1750 400
rect -1505 -100 -1405 400
rect -1325 -100 -1225 400
rect -1000 -100 -800 400
rect -600 -100 -400 400
rect -200 -100 0 400
rect 200 -100 400 400
rect 600 -100 800 400
rect 1000 -100 1200 400
rect 1400 -100 1600 400
rect 1800 -100 2000 400
rect 2200 -100 2400 400
rect 2600 -100 2800 400
rect 3000 -100 3200 400
rect 3400 -100 3600 400
rect 3800 -100 4000 400
rect 4200 -100 4400 400
rect 4550 -100 4750 400
<< pdiff >>
rect -3750 380 -3550 400
rect -3750 30 -3690 380
rect -3590 30 -3550 380
rect -3750 -100 -3550 30
rect -3350 380 -3150 400
rect -3350 30 -3300 380
rect -3200 30 -3150 380
rect -3350 -100 -3150 30
rect -2950 380 -2700 400
rect -2950 40 -2830 380
rect -2770 40 -2700 380
rect -2950 -100 -2700 40
rect -2600 340 -2400 400
rect -2600 30 -2540 340
rect -2460 30 -2400 340
rect -2600 -100 -2400 30
rect -2300 380 -2100 400
rect -2300 30 -2230 380
rect -2170 30 -2100 380
rect -2300 -100 -2100 30
rect -2000 380 -1850 400
rect -2000 40 -1960 380
rect -1890 40 -1850 380
rect -2000 -100 -1850 40
rect -1750 230 -1505 400
rect -1750 -60 -1680 230
rect -1620 -60 -1505 230
rect -1750 -100 -1505 -60
rect -1405 -100 -1325 400
rect -1225 290 -1000 400
rect -1225 40 -1120 290
rect -1080 40 -1000 290
rect -1225 -100 -1000 40
rect -800 270 -600 400
rect -800 30 -720 270
rect -680 30 -600 270
rect -800 -100 -600 30
rect -400 290 -200 400
rect -400 40 -320 290
rect -280 40 -200 290
rect -400 -100 -200 40
rect 0 270 200 400
rect 0 30 80 270
rect 120 30 200 270
rect 0 -100 200 30
rect 400 290 600 400
rect 400 40 480 290
rect 520 40 600 290
rect 400 -100 600 40
rect 800 270 1000 400
rect 800 30 880 270
rect 920 30 1000 270
rect 800 -100 1000 30
rect 1200 290 1400 400
rect 1200 40 1280 290
rect 1320 40 1400 290
rect 1200 -100 1400 40
rect 1600 270 1800 400
rect 1600 30 1680 270
rect 1720 30 1800 270
rect 1600 -100 1800 30
rect 2000 290 2200 400
rect 2000 40 2080 290
rect 2120 40 2200 290
rect 2000 -100 2200 40
rect 2400 270 2600 400
rect 2400 30 2480 270
rect 2520 30 2600 270
rect 2400 -100 2600 30
rect 2800 290 3000 400
rect 2800 40 2880 290
rect 2920 40 3000 290
rect 2800 -100 3000 40
rect 3200 270 3400 400
rect 3200 30 3280 270
rect 3320 30 3400 270
rect 3200 -100 3400 30
rect 3600 290 3800 400
rect 3600 40 3680 290
rect 3720 40 3800 290
rect 3600 -100 3800 40
rect 4000 380 4200 400
rect 4000 30 4050 380
rect 4150 30 4200 380
rect 4000 -100 4200 30
rect 4400 380 4550 400
rect 4400 40 4430 380
rect 4520 40 4550 380
rect 4400 -100 4550 40
rect 4750 380 4900 400
rect 4750 40 4780 380
rect 4870 40 4900 380
rect 4750 -100 4900 40
<< pdiffc >>
rect -3690 30 -3590 380
rect -3300 30 -3200 380
rect -2830 40 -2770 380
rect -2540 30 -2460 340
rect -2230 30 -2170 380
rect -1960 40 -1890 380
rect -1680 -60 -1620 230
rect -1120 40 -1080 290
rect -720 30 -680 270
rect -320 40 -280 290
rect 80 30 120 270
rect 480 40 520 290
rect 880 30 920 270
rect 1280 40 1320 290
rect 1680 30 1720 270
rect 2080 40 2120 290
rect 2480 30 2520 270
rect 2880 40 2920 290
rect 3280 30 3320 270
rect 3680 40 3720 290
rect 4050 30 4150 380
rect 4430 40 4520 380
rect 4780 40 4870 380
<< nsubdiff >>
rect -4040 1090 5120 1110
rect -4040 980 -3920 1090
rect -2270 980 -1970 1090
rect -320 980 310 1090
rect 1960 980 3350 1090
rect 5000 980 5120 1090
rect -4040 950 5120 980
rect -4040 910 -3850 950
rect -4040 -650 -4010 910
rect -3880 -600 -3850 910
rect 4980 940 5120 950
rect 4980 -590 5000 940
rect 5100 -590 5120 940
rect 4980 -600 5120 -590
rect -3880 -630 5120 -600
rect -3880 -650 -3840 -630
rect -4040 -740 -3840 -650
rect 1080 -730 1270 -630
rect 4990 -730 5120 -630
rect 1080 -740 5120 -730
rect -4040 -780 5120 -740
<< nsubdiffcont >>
rect -3920 980 -2270 1090
rect -1970 980 -320 1090
rect 310 980 1960 1090
rect 3350 980 5000 1090
rect -4010 -650 -3880 910
rect 5000 -590 5100 940
rect -3840 -740 1080 -630
rect 1270 -730 4990 -630
<< poly >>
rect -3550 590 -3350 600
rect -3550 510 -3540 590
rect -3360 510 -3350 590
rect -3550 400 -3350 510
rect -3150 590 -2950 600
rect -3150 510 -3140 590
rect -2960 510 -2950 590
rect -3150 400 -2950 510
rect -1505 590 -1405 600
rect -1505 510 -1495 590
rect -1415 510 -1405 590
rect -2700 400 -2600 500
rect -2400 400 -2300 500
rect -2100 490 -1750 500
rect -2100 430 -1980 490
rect -1870 430 -1750 490
rect -2100 420 -1750 430
rect -2100 400 -2000 420
rect -1850 400 -1750 420
rect -1505 400 -1405 510
rect -1325 591 -1225 600
rect -1325 511 -1315 591
rect -1235 511 -1225 591
rect -1325 400 -1225 511
rect -1000 580 -800 600
rect -1000 520 -980 580
rect -820 520 -800 580
rect -1000 400 -800 520
rect -600 580 -400 600
rect -600 520 -580 580
rect -420 520 -400 580
rect -600 400 -400 520
rect -200 580 0 600
rect -200 520 -180 580
rect -20 520 0 580
rect -200 400 0 520
rect 200 580 400 600
rect 200 520 220 580
rect 380 520 400 580
rect 200 400 400 520
rect 600 580 800 600
rect 600 520 620 580
rect 780 520 800 580
rect 600 400 800 520
rect 1000 580 1200 600
rect 1000 520 1020 580
rect 1180 520 1200 580
rect 1000 400 1200 520
rect 1400 580 1600 600
rect 1400 520 1420 580
rect 1580 520 1600 580
rect 1400 400 1600 520
rect 1800 580 2000 600
rect 1800 520 1820 580
rect 1980 520 2000 580
rect 1800 400 2000 520
rect 2200 580 2400 600
rect 2200 520 2220 580
rect 2380 520 2400 580
rect 2200 400 2400 520
rect 2600 580 2800 600
rect 2600 520 2620 580
rect 2780 520 2800 580
rect 2600 400 2800 520
rect 3000 580 3200 600
rect 3000 520 3020 580
rect 3180 520 3200 580
rect 3000 400 3200 520
rect 3400 580 3600 600
rect 3400 520 3420 580
rect 3580 520 3600 580
rect 3400 400 3600 520
rect 3800 590 4000 600
rect 3800 510 3810 590
rect 3990 510 4000 590
rect 3800 400 4000 510
rect 4200 590 4400 600
rect 4200 510 4210 590
rect 4390 510 4400 590
rect 4200 400 4400 510
rect 4550 590 4750 600
rect 4550 510 4560 590
rect 4740 510 4750 590
rect 4550 400 4750 510
rect -3550 -200 -3350 -100
rect -3150 -200 -2950 -100
rect -2700 -220 -2600 -100
rect -2700 -280 -2680 -220
rect -2620 -280 -2600 -220
rect -2700 -300 -2600 -280
rect -2400 -220 -2300 -100
rect -2100 -200 -2000 -100
rect -1850 -200 -1750 -100
rect -1505 -200 -1405 -100
rect -1325 -200 -1225 -100
rect -1000 -200 -800 -100
rect -600 -200 -400 -100
rect -200 -200 0 -100
rect 200 -200 400 -100
rect 600 -200 800 -100
rect 1000 -200 1200 -100
rect 1400 -200 1600 -100
rect 1800 -200 2000 -100
rect 2200 -200 2400 -100
rect 2600 -200 2800 -100
rect 3000 -200 3200 -100
rect 3400 -200 3600 -100
rect 3800 -200 4000 -100
rect 4200 -200 4400 -100
rect 4550 -200 4750 -100
rect -2400 -280 -2380 -220
rect -2320 -280 -2300 -220
rect -2400 -300 -2300 -280
<< polycont >>
rect -3540 510 -3360 590
rect -3140 510 -2960 590
rect -1495 510 -1415 590
rect -1980 430 -1870 490
rect -1315 511 -1235 591
rect -980 520 -820 580
rect -580 520 -420 580
rect -180 520 -20 580
rect 220 520 380 580
rect 620 520 780 580
rect 1020 520 1180 580
rect 1420 520 1580 580
rect 1820 520 1980 580
rect 2220 520 2380 580
rect 2620 520 2780 580
rect 3020 520 3180 580
rect 3420 520 3580 580
rect 3810 510 3990 590
rect 4210 510 4390 590
rect 4560 510 4740 590
rect -2680 -280 -2620 -220
rect -2380 -280 -2320 -220
<< locali >>
rect -4030 1090 5110 1100
rect -4030 980 -3920 1090
rect -2270 980 -1970 1090
rect -320 980 310 1090
rect 1960 980 3350 1090
rect 5000 980 5110 1090
rect -4030 960 5110 980
rect -4030 910 -3860 960
rect 4990 940 5110 960
rect -4030 -650 -4010 910
rect -3880 -610 -3860 910
rect 3450 920 4880 930
rect 3450 860 3460 920
rect 3540 860 4690 920
rect 4870 860 4880 920
rect 3450 850 4880 860
rect -3330 790 4880 800
rect -3330 730 -1980 790
rect -1870 780 -350 790
rect -1870 730 -1140 780
rect -3330 720 -1140 730
rect -1060 720 -350 780
rect -3330 600 -3180 720
rect -1160 710 -350 720
rect -250 710 450 790
rect 550 710 1250 790
rect 1350 710 2050 790
rect 2150 710 2850 790
rect 2950 710 3650 790
rect 3750 710 4690 790
rect 4870 710 4880 790
rect -1160 700 4880 710
rect -2850 610 -1450 690
rect -3710 590 -2950 600
rect -3710 510 -3540 590
rect -3360 510 -3140 590
rect -2960 510 -2950 590
rect -3710 500 -2950 510
rect -3710 380 -3570 500
rect -3710 30 -3690 380
rect -3590 30 -3570 380
rect -3710 -10 -3570 30
rect -3320 380 -3180 500
rect -3320 30 -3300 380
rect -3200 30 -3180 380
rect -3320 0 -3180 30
rect -2850 380 -2750 610
rect -2850 40 -2830 380
rect -2770 40 -2750 380
rect -2250 380 -2150 610
rect -1550 600 -1450 610
rect 4200 600 4400 700
rect -1550 591 3600 600
rect -1550 590 -1315 591
rect -1550 510 -1495 590
rect -1415 511 -1315 590
rect -1235 580 3600 591
rect -1235 520 -980 580
rect -820 520 -580 580
rect -420 520 -180 580
rect -20 520 220 580
rect 380 520 620 580
rect 780 520 1020 580
rect 1180 520 1420 580
rect 1580 520 1820 580
rect 1980 520 2220 580
rect 2380 520 2620 580
rect 2780 520 3020 580
rect 3180 520 3420 580
rect 3580 520 3600 580
rect -1235 511 3600 520
rect -1415 510 3600 511
rect -1550 500 3600 510
rect 3800 590 4880 600
rect 3800 510 3810 590
rect 3990 510 4210 590
rect 4390 510 4560 590
rect 4740 510 4880 590
rect 3800 500 4880 510
rect -2000 490 -1850 500
rect -2000 430 -1980 490
rect -1870 430 -1850 490
rect -2000 420 -1850 430
rect -2850 0 -2750 40
rect -2550 340 -2450 350
rect -2550 30 -2540 340
rect -2460 30 -2450 340
rect -2550 20 -2450 30
rect -2250 30 -2230 380
rect -2170 30 -2150 380
rect -2250 0 -2150 30
rect -1980 380 -1870 420
rect -1980 40 -1960 380
rect -1890 40 -1870 380
rect -1140 290 -1060 310
rect -340 290 -260 310
rect 460 290 540 310
rect -1140 270 -1120 290
rect -1080 270 -1060 290
rect -1980 0 -1870 40
rect -1700 230 -1600 250
rect -1700 -60 -1680 230
rect -1620 -60 -1600 230
rect -1140 60 -1130 270
rect -1070 60 -1060 270
rect -1140 40 -1120 60
rect -1080 40 -1060 60
rect -1140 20 -1060 40
rect -740 270 -660 290
rect -740 250 -720 270
rect -680 250 -660 270
rect -740 30 -720 40
rect -680 30 -660 40
rect -740 0 -660 30
rect -340 270 -320 290
rect -280 270 -260 290
rect -340 60 -330 270
rect -270 60 -260 270
rect -340 40 -320 60
rect -280 40 -260 60
rect -340 20 -260 40
rect 60 270 140 290
rect 60 250 80 270
rect 120 250 140 270
rect 60 30 80 50
rect 120 30 140 50
rect 60 0 140 30
rect 460 270 480 290
rect 520 270 540 290
rect 460 60 470 270
rect 530 60 540 270
rect 460 40 480 60
rect 520 40 540 60
rect 460 20 540 40
rect 860 270 940 500
rect 860 30 880 270
rect 920 30 940 270
rect 860 0 940 30
rect 1260 290 1340 310
rect 1260 270 1280 290
rect 1320 270 1340 290
rect 1260 60 1270 270
rect 1330 60 1340 270
rect 1260 40 1280 60
rect 1320 40 1340 60
rect 1260 20 1340 40
rect 1660 270 1740 500
rect 4040 380 4160 500
rect 1660 30 1680 270
rect 1720 30 1740 270
rect 1660 0 1740 30
rect 2060 290 2140 310
rect 2860 290 2940 310
rect 3660 290 3740 310
rect 2060 270 2080 290
rect 2120 270 2140 290
rect 2060 60 2070 270
rect 2130 60 2140 270
rect 2060 40 2080 60
rect 2120 40 2140 60
rect 2060 20 2140 40
rect 2460 270 2540 290
rect 2460 250 2480 270
rect 2520 250 2540 270
rect 2460 30 2480 40
rect 2520 30 2540 40
rect 2460 0 2540 30
rect 2860 270 2880 290
rect 2920 270 2940 290
rect 2860 60 2870 270
rect 2930 60 2940 270
rect 2860 40 2880 60
rect 2920 40 2940 60
rect 2860 20 2940 40
rect 3260 270 3340 290
rect 3260 250 3280 270
rect 3320 250 3340 270
rect 3260 30 3280 40
rect 3320 30 3340 40
rect 3260 0 3340 30
rect 3660 270 3680 290
rect 3720 270 3740 290
rect 3660 60 3670 270
rect 3730 60 3740 270
rect 3660 40 3680 60
rect 3720 40 3740 60
rect 3660 20 3740 40
rect 4040 30 4050 380
rect 4150 30 4160 380
rect 4040 0 4160 30
rect 4420 380 4530 500
rect 4420 40 4430 380
rect 4520 40 4530 380
rect 4420 10 4530 40
rect 4770 380 4880 500
rect 4770 40 4780 380
rect 4870 40 4880 380
rect 4770 10 4880 40
rect -1700 -200 -1600 -60
rect -2700 -220 -1600 -200
rect -2700 -280 -2680 -220
rect -2620 -280 -2380 -220
rect -2320 -280 -1600 -220
rect -2700 -300 -1600 -280
rect -2550 -330 4670 -320
rect -2550 -410 -2540 -330
rect -2460 -400 50 -330
rect 150 -400 2450 -330
rect -2460 -410 2450 -400
rect 2550 -410 4450 -330
rect 4660 -410 4670 -330
rect -2550 -420 4670 -410
rect -1130 -470 4670 -460
rect -1130 -550 -750 -470
rect -650 -550 3250 -470
rect 3350 -550 4450 -470
rect 4660 -550 4670 -470
rect -1130 -560 4670 -550
rect 4990 -590 5000 940
rect 5100 -590 5110 940
rect 4990 -610 5110 -590
rect -3880 -630 5110 -610
rect -3880 -650 -3840 -630
rect -4030 -740 -3840 -650
rect 1080 -730 1270 -630
rect 4990 -730 5110 -630
rect 1080 -740 5110 -730
rect -4030 -770 5110 -740
<< viali >>
rect 3460 860 3540 920
rect 4690 860 4870 920
rect -1980 730 -1870 790
rect -1140 720 -1060 780
rect -350 710 -250 790
rect 450 710 550 790
rect 1250 710 1350 790
rect 2050 710 2150 790
rect 2850 710 2950 790
rect 3650 710 3750 790
rect 4690 710 4870 790
rect 3460 520 3540 580
rect -1970 430 -1880 490
rect -2540 70 -2460 300
rect -1680 -30 -1620 200
rect -1130 60 -1120 270
rect -1120 60 -1080 270
rect -1080 60 -1070 270
rect -740 40 -720 250
rect -720 40 -680 250
rect -680 40 -660 250
rect -330 60 -320 270
rect -320 60 -280 270
rect -280 60 -270 270
rect 60 50 80 250
rect 80 50 120 250
rect 120 50 140 250
rect 470 60 480 270
rect 480 60 520 270
rect 520 60 530 270
rect 1270 60 1280 270
rect 1280 60 1320 270
rect 1320 60 1330 270
rect 2070 60 2080 270
rect 2080 60 2120 270
rect 2120 60 2130 270
rect 2460 40 2480 250
rect 2480 40 2520 250
rect 2520 40 2540 250
rect 2870 60 2880 270
rect 2880 60 2920 270
rect 2920 60 2930 270
rect 3260 40 3280 250
rect 3280 40 3320 250
rect 3320 40 3340 250
rect 3670 60 3680 270
rect 3680 60 3720 270
rect 3720 60 3730 270
rect -2540 -410 -2460 -330
rect 50 -400 150 -330
rect 2450 -410 2550 -330
rect 4450 -410 4660 -330
rect -750 -550 -650 -470
rect 3250 -550 3350 -470
rect 4450 -550 4660 -470
<< metal1 >>
rect 3450 920 3550 930
rect 3450 860 3460 920
rect 3540 860 3550 920
rect -1990 790 -1860 800
rect -1990 730 -1980 790
rect -1870 730 -1860 790
rect -1990 490 -1860 730
rect -1990 430 -1970 490
rect -1880 430 -1860 490
rect -1990 420 -1860 430
rect -1160 780 -1040 800
rect -1160 720 -1140 780
rect -1060 720 -1040 780
rect -2550 300 -2450 350
rect -2550 70 -2540 300
rect -2460 70 -2450 300
rect -1160 270 -1040 720
rect -360 790 -240 800
rect -360 710 -350 790
rect -250 710 -240 790
rect -2550 -330 -2450 70
rect -2550 -410 -2540 -330
rect -2460 -410 -2450 -330
rect -2550 -420 -2450 -410
rect -1700 200 -1600 250
rect -1700 -30 -1680 200
rect -1620 -30 -1600 200
rect -1160 60 -1130 270
rect -1070 60 -1040 270
rect -1160 0 -1040 60
rect -760 250 -640 320
rect -760 40 -740 250
rect -660 40 -640 250
rect -1700 -930 -1600 -30
rect -760 -470 -640 40
rect -360 270 -240 710
rect 440 790 560 800
rect 440 710 450 790
rect 550 710 560 790
rect -360 60 -330 270
rect -270 60 -240 270
rect -360 0 -240 60
rect 40 250 160 330
rect 40 50 60 250
rect 140 50 160 250
rect 40 -330 160 50
rect 440 270 560 710
rect 440 60 470 270
rect 530 60 560 270
rect 440 0 560 60
rect 1240 790 1360 800
rect 1240 710 1250 790
rect 1350 710 1360 790
rect 1240 270 1360 710
rect 1240 60 1270 270
rect 1330 60 1360 270
rect 1240 0 1360 60
rect 2040 790 2160 800
rect 2040 710 2050 790
rect 2150 710 2160 790
rect 2040 270 2160 710
rect 2840 790 2960 800
rect 2840 710 2850 790
rect 2950 710 2960 790
rect 2040 60 2070 270
rect 2130 60 2160 270
rect 2040 0 2160 60
rect 2440 250 2560 330
rect 2440 40 2460 250
rect 2540 40 2560 250
rect 40 -400 50 -330
rect 150 -400 160 -330
rect 40 -420 160 -400
rect 2440 -330 2560 40
rect 2840 270 2960 710
rect 3450 580 3550 860
rect 4680 920 5310 930
rect 4680 860 4690 920
rect 4870 860 5310 920
rect 4680 850 5310 860
rect 3450 520 3460 580
rect 3540 520 3550 580
rect 3450 500 3550 520
rect 3640 790 3760 800
rect 3640 710 3650 790
rect 3750 710 3760 790
rect 2840 60 2870 270
rect 2930 60 2960 270
rect 2840 0 2960 60
rect 3240 250 3360 320
rect 3240 40 3260 250
rect 3340 40 3360 250
rect 2440 -410 2450 -330
rect 2550 -410 2560 -330
rect 2440 -420 2560 -410
rect -760 -550 -750 -470
rect -650 -550 -640 -470
rect -760 -560 -640 -550
rect 3240 -470 3360 40
rect 3640 270 3760 710
rect 4680 790 5310 800
rect 4680 710 4690 790
rect 4870 710 5310 790
rect 4680 700 5310 710
rect 3640 60 3670 270
rect 3730 60 3760 270
rect 3640 0 3760 60
rect 4440 -330 5470 -320
rect 4440 -410 4450 -330
rect 4660 -410 5470 -330
rect 4440 -420 5470 -410
rect 3240 -550 3250 -470
rect 3350 -550 3360 -470
rect 3240 -560 3360 -550
rect 4440 -470 5470 -460
rect 4440 -550 4450 -470
rect 4660 -550 5470 -470
rect 4440 -560 5470 -550
<< end >>
