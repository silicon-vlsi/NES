magic
tech sky130A
timestamp 1767954981
<< nwell >>
rect -20 135 310 315
<< nmos >>
rect 75 51 90 93
rect 120 51 135 93
rect 165 51 180 93
rect 210 51 225 93
<< pmos >>
rect 45 160 60 219
rect 90 160 105 219
rect 190 160 205 219
rect 235 160 250 219
<< ndiff >>
rect 48 79 75 93
rect 48 62 52 79
rect 69 62 75 79
rect 48 51 75 62
rect 90 79 120 93
rect 90 62 96 79
rect 114 62 120 79
rect 90 51 120 62
rect 135 79 165 93
rect 135 62 141 79
rect 159 62 165 79
rect 135 51 165 62
rect 180 79 210 93
rect 180 62 186 79
rect 204 62 210 79
rect 180 51 210 62
rect 225 79 253 93
rect 225 62 231 79
rect 249 62 253 79
rect 225 51 253 62
<< pdiff >>
rect 18 211 45 219
rect 18 194 22 211
rect 39 194 45 211
rect 18 160 45 194
rect 60 211 90 219
rect 60 194 66 211
rect 84 194 90 211
rect 60 160 90 194
rect 105 211 133 219
rect 105 194 111 211
rect 129 194 133 211
rect 105 160 133 194
rect 163 211 190 219
rect 163 194 167 211
rect 184 194 190 211
rect 163 160 190 194
rect 205 211 235 219
rect 205 194 211 211
rect 229 194 235 211
rect 205 160 235 194
rect 250 211 278 219
rect 250 194 256 211
rect 274 194 278 211
rect 250 160 278 194
<< ndiffc >>
rect 52 62 69 79
rect 96 62 114 79
rect 141 62 159 79
rect 186 62 204 79
rect 231 62 249 79
<< pdiffc >>
rect 22 194 39 211
rect 66 194 84 211
rect 111 194 129 211
rect 167 194 184 211
rect 211 194 229 211
rect 256 194 274 211
<< psubdiff >>
rect 30 7 264 24
rect 30 -10 45 7
rect 62 -10 95 7
rect 114 -10 140 7
rect 159 -10 185 7
rect 204 -10 231 7
rect 249 -10 264 7
rect 30 -24 264 -10
<< nsubdiff >>
rect 0 278 291 295
rect 0 261 15 278
rect 32 261 65 278
rect 84 261 111 278
rect 129 261 160 278
rect 177 261 210 278
rect 229 261 256 278
rect 274 261 291 278
rect 0 246 291 261
<< psubdiffcont >>
rect 45 -10 62 7
rect 95 -10 114 7
rect 140 -10 159 7
rect 185 -10 204 7
rect 231 -10 249 7
<< nsubdiffcont >>
rect 15 261 32 278
rect 65 261 84 278
rect 111 261 129 278
rect 160 261 177 278
rect 210 261 229 278
rect 256 261 274 278
<< poly >>
rect 45 219 60 232
rect 90 219 105 232
rect 190 219 205 232
rect 235 219 250 232
rect 45 143 60 160
rect 15 135 60 143
rect 15 118 20 135
rect 37 125 60 135
rect 90 125 105 160
rect 190 125 205 160
rect 235 143 250 160
rect 235 135 280 143
rect 235 125 255 135
rect 37 118 135 125
rect 15 110 135 118
rect 75 93 90 110
rect 120 93 135 110
rect 165 118 255 125
rect 272 118 280 135
rect 165 110 280 118
rect 165 93 180 110
rect 210 93 225 110
rect 75 38 90 51
rect 120 38 135 51
rect 165 38 180 51
rect 210 38 225 51
<< polycont >>
rect 20 118 37 135
rect 255 118 272 135
<< locali >>
rect 0 278 291 295
rect 0 261 15 278
rect 32 261 65 278
rect 84 261 111 278
rect 129 261 160 278
rect 177 261 210 278
rect 229 261 256 278
rect 274 261 291 278
rect 0 246 291 261
rect 17 219 42 246
rect 60 223 88 228
rect 17 211 43 219
rect 17 200 22 211
rect 18 194 22 200
rect 39 194 43 211
rect 60 201 66 223
rect 18 160 43 194
rect 62 194 66 201
rect 84 194 88 223
rect 108 219 133 246
rect 62 159 88 194
rect 107 211 133 219
rect 107 194 111 211
rect 129 194 133 211
rect 107 159 133 194
rect 163 223 188 228
rect 163 194 167 223
rect 185 206 188 223
rect 252 223 278 228
rect 184 194 188 206
rect 163 160 188 194
rect 207 211 233 219
rect 207 194 211 211
rect 229 194 233 211
rect 207 182 233 194
rect 207 165 211 182
rect 229 165 233 182
rect 207 159 233 165
rect 252 206 254 223
rect 272 211 278 223
rect 252 194 256 206
rect 274 194 278 211
rect 252 160 278 194
rect 15 135 45 143
rect 15 118 20 135
rect 37 118 45 135
rect 15 110 45 118
rect 250 135 280 143
rect 250 118 255 135
rect 272 118 280 135
rect 250 110 280 118
rect 48 79 73 93
rect 48 62 52 79
rect 69 62 73 79
rect 48 24 73 62
rect 92 81 118 93
rect 92 62 96 81
rect 114 62 118 81
rect 92 51 118 62
rect 137 79 163 93
rect 137 62 141 79
rect 159 62 163 79
rect 137 51 163 62
rect 182 81 208 93
rect 182 62 186 81
rect 204 62 208 81
rect 182 51 208 62
rect 227 79 253 93
rect 227 62 231 79
rect 249 62 253 79
rect 227 51 253 62
rect 138 24 163 51
rect 228 24 253 51
rect 30 7 264 24
rect 30 -10 45 7
rect 62 -10 95 7
rect 114 -10 140 7
rect 159 -10 185 7
rect 204 -10 231 7
rect 249 -10 264 7
rect 30 -25 264 -10
<< viali >>
rect 15 261 32 278
rect 65 261 84 278
rect 111 261 129 278
rect 160 261 177 278
rect 210 261 229 278
rect 256 261 274 278
rect 66 211 84 223
rect 66 206 84 211
rect 167 211 185 223
rect 167 206 184 211
rect 184 206 185 211
rect 211 165 229 182
rect 254 211 272 223
rect 254 206 256 211
rect 256 206 272 211
rect 20 118 37 135
rect 255 118 272 135
rect 96 79 114 81
rect 96 64 114 79
rect 186 79 204 81
rect 186 64 204 79
rect 45 -10 62 7
rect 95 -10 114 7
rect 140 -10 159 7
rect 185 -10 204 7
rect 231 -10 249 7
<< metal1 >>
rect 0 278 291 295
rect 0 261 15 278
rect 32 261 65 278
rect 84 261 111 278
rect 129 261 160 278
rect 177 261 210 278
rect 229 261 256 278
rect 274 261 291 278
rect 0 246 291 261
rect 60 223 278 228
rect 60 206 66 223
rect 84 206 167 223
rect 185 206 254 223
rect 272 206 278 223
rect 60 201 278 206
rect 62 200 278 201
rect 204 182 235 186
rect 204 165 211 182
rect 229 165 235 182
rect 204 160 235 165
rect 15 142 45 143
rect 15 135 46 142
rect 15 118 20 135
rect 37 118 46 135
rect 15 111 46 118
rect 15 110 45 111
rect 207 86 233 160
rect 250 135 280 143
rect 250 118 255 135
rect 272 118 280 135
rect 250 110 280 118
rect 90 81 233 86
rect 90 64 96 81
rect 114 64 186 81
rect 204 64 233 81
rect 90 60 233 64
rect 30 7 264 24
rect 30 -10 45 7
rect 62 -10 95 7
rect 114 -10 140 7
rect 159 -10 185 7
rect 204 -10 231 7
rect 249 -10 264 7
rect 30 -25 264 -10
<< end >>
