magic
tech sky130A
timestamp 1767943905
<< fence >>
rect 0 0 480 270
<< nwell >>
rect -20 135 505 315
<< nmos >>
rect 45 51 60 93
rect 90 51 105 93
rect 135 51 150 93
rect 180 51 195 93
rect 290 51 305 93
rect 335 51 350 93
rect 380 51 395 93
rect 425 51 440 93
<< pmos >>
rect 75 160 90 219
rect 120 160 135 219
rect 165 160 180 219
rect 210 160 225 219
rect 255 160 270 219
rect 300 160 315 219
rect 345 160 360 219
rect 390 160 405 219
<< ndiff >>
rect 18 79 45 93
rect 18 62 22 79
rect 39 62 45 79
rect 18 51 45 62
rect 60 89 90 93
rect 60 72 67 89
rect 84 72 90 89
rect 60 51 90 72
rect 105 83 135 93
rect 105 66 112 83
rect 129 66 135 83
rect 105 51 135 66
rect 150 89 180 93
rect 150 72 157 89
rect 174 72 180 89
rect 150 51 180 72
rect 195 82 225 93
rect 195 65 203 82
rect 220 65 225 82
rect 195 51 225 65
rect 263 79 290 93
rect 263 62 267 79
rect 284 62 290 79
rect 263 51 290 62
rect 305 79 335 93
rect 305 62 311 79
rect 329 62 335 79
rect 305 51 335 62
rect 350 79 380 93
rect 350 62 356 79
rect 374 62 380 79
rect 350 51 380 62
rect 395 79 425 93
rect 395 62 401 79
rect 419 62 425 79
rect 395 51 425 62
rect 440 79 470 93
rect 440 62 446 79
rect 464 62 470 79
rect 440 51 470 62
<< pdiff >>
rect 48 211 75 219
rect 48 194 52 211
rect 69 194 75 211
rect 48 160 75 194
rect 90 211 120 219
rect 90 194 96 211
rect 114 194 120 211
rect 90 160 120 194
rect 135 211 165 219
rect 135 194 141 211
rect 159 194 165 211
rect 135 160 165 194
rect 180 211 210 219
rect 180 194 186 211
rect 204 194 210 211
rect 180 160 210 194
rect 225 211 255 219
rect 225 194 231 211
rect 249 194 255 211
rect 225 160 255 194
rect 270 211 300 219
rect 270 194 276 211
rect 294 194 300 211
rect 270 160 300 194
rect 315 211 345 219
rect 315 194 321 211
rect 339 194 345 211
rect 315 160 345 194
rect 360 211 390 219
rect 360 194 366 211
rect 384 194 390 211
rect 360 160 390 194
rect 405 211 432 219
rect 405 194 411 211
rect 428 194 432 211
rect 405 160 432 194
<< ndiffc >>
rect 22 62 39 79
rect 67 72 84 89
rect 112 66 129 83
rect 157 72 174 89
rect 203 65 220 82
rect 267 62 284 79
rect 311 62 329 79
rect 356 62 374 79
rect 401 62 419 79
rect 446 62 464 79
<< pdiffc >>
rect 52 194 69 211
rect 96 194 114 211
rect 141 194 159 211
rect 186 194 204 211
rect 231 194 249 211
rect 276 194 294 211
rect 321 194 339 211
rect 366 194 384 211
rect 411 194 428 211
<< psubdiff >>
rect 0 7 479 24
rect 0 -10 15 7
rect 32 -10 60 7
rect 80 -10 105 7
rect 125 -10 150 7
rect 170 -10 201 7
rect 219 -10 260 7
rect 277 -10 305 7
rect 325 -10 350 7
rect 370 -10 395 7
rect 415 -10 446 7
rect 464 -10 479 7
rect 0 -24 479 -10
rect 225 -25 255 -24
<< nsubdiff >>
rect 441 295 480 296
rect 0 278 480 295
rect 0 261 45 278
rect 62 261 90 278
rect 110 261 135 278
rect 155 261 180 278
rect 200 261 225 278
rect 245 261 270 278
rect 290 261 315 278
rect 335 261 360 278
rect 380 261 411 278
rect 429 261 480 278
rect 0 246 480 261
<< psubdiffcont >>
rect 15 -10 32 7
rect 60 -10 80 7
rect 105 -10 125 7
rect 150 -10 170 7
rect 201 -10 219 7
rect 260 -10 277 7
rect 305 -10 325 7
rect 350 -10 370 7
rect 395 -10 415 7
rect 446 -10 464 7
<< nsubdiffcont >>
rect 45 261 62 278
rect 90 261 110 278
rect 135 261 155 278
rect 180 261 200 278
rect 225 261 245 278
rect 270 261 290 278
rect 315 261 335 278
rect 360 261 380 278
rect 411 261 429 278
<< poly >>
rect 75 219 90 232
rect 120 219 135 232
rect 165 219 180 232
rect 210 219 225 232
rect 255 219 270 232
rect 300 219 315 232
rect 345 219 360 232
rect 390 219 405 232
rect 75 125 90 160
rect 120 143 135 160
rect 165 143 180 160
rect 120 135 180 143
rect 120 125 140 135
rect 45 118 140 125
rect 157 125 180 135
rect 210 125 225 160
rect 157 118 225 125
rect 45 110 225 118
rect 255 125 270 160
rect 300 125 315 160
rect 345 125 360 160
rect 390 143 405 160
rect 390 135 440 143
rect 390 125 410 135
rect 255 118 410 125
rect 427 118 440 135
rect 255 110 440 118
rect 45 93 60 110
rect 90 93 105 110
rect 135 93 150 110
rect 180 93 195 110
rect 290 93 305 110
rect 335 93 350 110
rect 380 93 395 110
rect 425 93 440 110
rect 45 38 60 51
rect 90 38 105 51
rect 135 38 150 51
rect 180 38 195 51
rect 290 38 305 51
rect 335 38 350 51
rect 380 38 395 51
rect 425 38 440 51
<< polycont >>
rect 140 118 157 135
rect 410 118 427 135
<< locali >>
rect 441 295 480 296
rect 0 278 480 295
rect 0 261 45 278
rect 62 261 90 278
rect 110 261 135 278
rect 155 261 180 278
rect 200 261 225 278
rect 245 261 270 278
rect 290 261 315 278
rect 335 261 360 278
rect 380 261 411 278
rect 429 261 480 278
rect 0 246 480 261
rect 48 211 73 246
rect 137 219 162 246
rect 227 219 252 246
rect 317 219 342 246
rect 48 194 52 211
rect 69 194 73 211
rect 48 160 73 194
rect 92 211 118 219
rect 92 187 96 211
rect 114 187 118 211
rect 92 160 118 187
rect 137 211 163 219
rect 137 194 141 211
rect 159 194 163 211
rect 137 160 163 194
rect 182 211 208 219
rect 182 188 186 211
rect 204 188 208 211
rect 182 160 208 188
rect 227 211 253 219
rect 227 194 231 211
rect 249 194 253 211
rect 227 160 253 194
rect 272 211 298 219
rect 272 188 276 211
rect 294 188 298 211
rect 272 160 298 188
rect 317 211 343 219
rect 317 194 321 211
rect 339 194 343 211
rect 317 160 343 194
rect 362 211 388 219
rect 362 194 366 211
rect 384 205 388 211
rect 362 188 367 194
rect 385 188 388 205
rect 362 160 388 188
rect 407 211 432 246
rect 407 194 411 211
rect 428 194 432 211
rect 407 160 432 194
rect 135 135 165 143
rect 135 118 140 135
rect 157 118 165 135
rect 135 110 165 118
rect 405 135 440 143
rect 405 118 410 135
rect 427 118 440 135
rect 405 110 440 118
rect 18 79 42 93
rect 18 62 22 79
rect 39 62 42 79
rect 59 89 92 93
rect 59 68 67 89
rect 84 68 92 89
rect 109 83 132 93
rect 18 50 42 62
rect 109 66 112 83
rect 129 66 132 83
rect 149 89 182 93
rect 149 68 157 89
rect 174 68 182 89
rect 199 82 225 93
rect 263 92 288 93
rect 109 50 132 66
rect 199 65 203 82
rect 220 65 225 82
rect 199 50 225 65
rect 18 32 225 50
rect 262 79 288 92
rect 262 62 267 79
rect 284 62 288 79
rect 262 14 288 62
rect 307 84 333 93
rect 307 79 313 84
rect 307 62 311 79
rect 330 67 333 84
rect 329 62 333 67
rect 307 51 333 62
rect 352 92 378 93
rect 352 79 379 92
rect 352 62 356 79
rect 374 62 379 79
rect 352 51 379 62
rect 397 84 423 93
rect 397 62 401 84
rect 418 79 423 84
rect 419 62 423 79
rect 397 51 423 62
rect 442 88 468 93
rect 442 79 469 88
rect 442 62 446 79
rect 464 62 469 79
rect 442 51 469 62
rect 353 34 379 51
rect 443 35 469 51
rect 353 14 380 34
rect 443 14 470 35
rect 0 7 479 14
rect 0 -10 15 7
rect 32 -10 60 7
rect 80 -10 105 7
rect 125 -10 150 7
rect 170 -10 201 7
rect 219 -10 260 7
rect 277 -10 305 7
rect 325 -10 350 7
rect 370 -10 395 7
rect 415 -10 446 7
rect 464 -10 479 7
rect 0 -25 479 -10
<< viali >>
rect 45 261 62 278
rect 90 261 110 278
rect 135 261 155 278
rect 180 261 200 278
rect 225 261 245 278
rect 270 261 290 278
rect 315 261 335 278
rect 360 261 380 278
rect 411 261 429 278
rect 96 194 114 204
rect 96 187 114 194
rect 186 194 204 205
rect 186 188 204 194
rect 276 194 294 205
rect 276 188 294 194
rect 367 194 384 205
rect 384 194 385 205
rect 367 188 385 194
rect 140 118 157 135
rect 410 118 427 135
rect 22 62 39 79
rect 67 72 84 84
rect 67 67 84 72
rect 157 72 174 84
rect 157 67 174 72
rect 313 79 330 84
rect 313 67 329 79
rect 329 67 330 79
rect 401 79 418 84
rect 401 67 418 79
rect 15 -10 32 7
rect 60 -10 80 7
rect 105 -10 125 7
rect 150 -10 170 7
rect 201 -10 219 7
rect 260 -10 277 7
rect 305 -10 325 7
rect 350 -10 370 7
rect 395 -10 415 7
rect 446 -10 464 7
<< metal1 >>
rect 441 295 480 296
rect 0 278 480 295
rect 0 261 45 278
rect 62 261 90 278
rect 110 261 135 278
rect 155 261 180 278
rect 200 261 225 278
rect 245 261 270 278
rect 290 261 315 278
rect 335 261 360 278
rect 380 261 411 278
rect 429 261 480 278
rect 0 246 480 261
rect 17 205 388 214
rect 17 204 186 205
rect 17 187 96 204
rect 114 188 186 204
rect 204 188 276 205
rect 294 188 367 205
rect 385 188 388 205
rect 114 187 388 188
rect 17 177 388 187
rect 18 79 44 177
rect 91 176 388 177
rect 135 142 165 143
rect 135 135 166 142
rect 135 118 140 135
rect 157 118 166 135
rect 135 111 166 118
rect 405 135 440 143
rect 405 118 410 135
rect 427 118 440 135
rect 135 110 165 111
rect 405 110 440 118
rect 18 62 22 79
rect 39 62 44 79
rect 18 51 44 62
rect 60 84 423 90
rect 60 67 67 84
rect 84 67 157 84
rect 174 67 313 84
rect 330 67 401 84
rect 418 67 423 84
rect 60 58 423 67
rect 0 7 479 24
rect 0 -10 15 7
rect 32 -10 60 7
rect 80 -10 105 7
rect 125 -10 150 7
rect 170 -10 201 7
rect 219 -10 260 7
rect 277 -10 305 7
rect 325 -10 350 7
rect 370 -10 395 7
rect 415 -10 446 7
rect 464 -10 479 7
rect 0 -25 479 -10
<< labels >>
rlabel nwell 15 251 465 287 1 vdd
port 1 n
rlabel metal1 12 -21 470 13 1 gnd
port 2 n
rlabel metal1 140 114 163 129 1 a
port 3 n
rlabel metal1 408 116 431 131 1 b
port 4 n
rlabel metal1 23 111 38 125 1 out
port 5 n
<< end >>
