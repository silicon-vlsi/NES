magic
tech sky130A
magscale 1 2
timestamp 1769684413
<< nwell >>
rect 2338 582 2564 584
rect 2278 260 2564 582
rect 2338 -378 2564 260
rect 2322 -700 2564 -378
<< locali >>
rect 998 527 2420 561
rect 954 -433 2420 -399
<< viali >>
rect 1566 356 1610 423
rect 2217 322 2258 445
rect 1168 216 1271 253
rect 1323 215 1377 249
rect 1833 218 1907 253
rect 1966 218 2024 252
rect 1321 -557 1378 -522
rect 987 -737 1046 -702
rect 1159 -739 1212 -703
rect 1447 -734 1514 -695
rect 1617 -738 1676 -701
rect 1817 -794 1851 -720
rect 1923 -794 1957 -720
rect 2084 -757 2118 -712
rect 2258 -748 2299 -625
<< metal1 >>
rect 838 580 2648 592
rect 838 505 2340 580
rect 2412 505 2648 580
rect 838 496 2648 505
rect 2205 445 2643 461
rect 1812 439 1921 441
rect 1559 424 1921 439
rect 1559 423 1612 424
rect 1559 356 1566 423
rect 1610 360 1612 423
rect 1690 360 1921 424
rect 1610 356 1921 360
rect 1559 344 1921 356
rect 1156 253 1283 261
rect 1156 216 1168 253
rect 1271 216 1283 253
rect 1156 199 1184 216
rect 1260 199 1283 216
rect 1156 193 1283 199
rect 1311 255 1394 261
rect 1311 202 1321 255
rect 1373 249 1394 255
rect 1377 215 1394 249
rect 1373 202 1394 215
rect 1812 253 1921 344
rect 2205 322 2217 445
rect 2258 322 2643 445
rect 2205 310 2643 322
rect 1812 218 1833 253
rect 1907 218 1921 253
rect 1812 215 1921 218
rect 1953 252 2049 263
rect 1953 246 1966 252
rect 2024 246 2049 252
rect 1812 212 1920 215
rect 1311 192 1394 202
rect 1953 193 1965 246
rect 2033 193 2049 246
rect 1953 187 2049 193
rect 2228 38 2561 48
rect 2228 -37 2481 38
rect 2553 -37 2561 38
rect 2228 -48 2561 -37
rect 845 -80 1181 -79
rect 845 -135 980 -80
rect 1064 -135 1181 -80
rect 1260 -135 2308 -79
rect 843 -173 2309 -169
rect 843 -176 1314 -173
rect 843 -232 1146 -176
rect 1217 -230 1314 -176
rect 1395 -230 2309 -173
rect 1217 -232 2309 -230
rect 843 -234 2309 -232
rect 845 -328 1441 -276
rect 1523 -278 2309 -276
rect 1523 -328 1963 -278
rect 845 -331 1963 -328
rect 2042 -331 2309 -278
rect 845 -332 2309 -331
rect 954 -378 2428 -368
rect 954 -453 2338 -378
rect 2410 -453 2428 -378
rect 954 -464 2428 -453
rect 1305 -522 1397 -508
rect 1305 -557 1321 -522
rect 1378 -557 1397 -522
rect 1305 -560 1397 -557
rect 975 -653 1070 -622
rect 975 -737 987 -653
rect 1046 -737 1070 -653
rect 975 -745 1070 -737
rect 1143 -656 1226 -623
rect 1305 -642 1321 -560
rect 1378 -642 1397 -560
rect 2247 -625 2685 -611
rect 1305 -643 1397 -642
rect 1143 -723 1151 -656
rect 1217 -723 1226 -656
rect 1143 -739 1159 -723
rect 1212 -739 1226 -723
rect 1143 -745 1226 -739
rect 1434 -647 1530 -625
rect 1434 -734 1447 -647
rect 1514 -734 1530 -647
rect 1434 -745 1530 -734
rect 1599 -664 1702 -653
rect 1599 -719 1614 -664
rect 1686 -719 1702 -664
rect 1599 -738 1617 -719
rect 1676 -738 1702 -719
rect 1599 -745 1702 -738
rect 1807 -720 1974 -695
rect 1807 -794 1817 -720
rect 1851 -794 1923 -720
rect 1957 -794 1974 -720
rect 1807 -808 1974 -794
rect 2062 -712 2145 -694
rect 2062 -739 2084 -712
rect 2118 -739 2145 -712
rect 2062 -792 2076 -739
rect 2129 -792 2145 -739
rect 2247 -748 2258 -625
rect 2299 -748 2685 -625
rect 2247 -762 2685 -748
rect 2062 -807 2145 -792
rect 819 -922 2641 -911
rect 819 -997 2481 -922
rect 2553 -997 2641 -922
rect 819 -1008 2641 -997
rect 2150 -1039 2467 -1038
rect 1009 -1053 2467 -1039
rect 1009 -1111 1314 -1053
rect 1385 -1055 2467 -1053
rect 1385 -1109 2077 -1055
rect 2129 -1109 2467 -1055
rect 1385 -1111 2467 -1109
rect 1009 -1124 2467 -1111
rect 2150 -1125 2467 -1124
<< via1 >>
rect 2340 505 2412 580
rect 1612 360 1690 424
rect 1184 216 1260 253
rect 1184 199 1260 216
rect 1321 249 1373 255
rect 1321 215 1323 249
rect 1323 215 1373 249
rect 1321 202 1373 215
rect 1965 218 1966 246
rect 1966 218 2024 246
rect 2024 218 2033 246
rect 1965 193 2033 218
rect 2481 -37 2553 38
rect 980 -135 1064 -80
rect 1181 -135 1260 -79
rect 1146 -232 1217 -176
rect 1314 -230 1395 -173
rect 1441 -328 1523 -276
rect 1963 -331 2042 -278
rect 2338 -453 2410 -378
rect 987 -702 1046 -653
rect 987 -706 1046 -702
rect 1321 -642 1378 -560
rect 1151 -703 1217 -656
rect 1151 -723 1159 -703
rect 1159 -723 1212 -703
rect 1212 -723 1217 -703
rect 1447 -695 1514 -647
rect 1447 -706 1514 -695
rect 1614 -701 1686 -664
rect 1614 -719 1617 -701
rect 1617 -719 1676 -701
rect 1676 -719 1686 -701
rect 2076 -757 2084 -739
rect 2084 -757 2118 -739
rect 2118 -757 2129 -739
rect 2076 -792 2129 -757
rect 2481 -997 2553 -922
rect 1314 -1111 1385 -1053
rect 2077 -1109 2129 -1055
<< metal2 >>
rect 2332 580 2420 591
rect 2332 505 2340 580
rect 2412 505 2420 580
rect 1599 424 1702 439
rect 1599 360 1612 424
rect 1690 360 1702 424
rect 1176 253 1267 261
rect 1176 199 1184 253
rect 1260 199 1267 253
rect 975 -80 1070 -71
rect 975 -135 980 -80
rect 1064 -135 1070 -80
rect 975 -653 1070 -135
rect 1176 -79 1267 199
rect 1176 -135 1181 -79
rect 1260 -135 1267 -79
rect 1176 -141 1267 -135
rect 1310 255 1401 262
rect 1310 202 1321 255
rect 1373 202 1401 255
rect 975 -706 987 -653
rect 1046 -706 1070 -653
rect 975 -745 1070 -706
rect 1143 -176 1226 -169
rect 1143 -232 1146 -176
rect 1217 -232 1226 -176
rect 1143 -656 1226 -232
rect 1310 -173 1401 202
rect 1310 -230 1314 -173
rect 1395 -230 1401 -173
rect 1310 -237 1401 -230
rect 1434 -328 1441 -276
rect 1523 -328 1530 -276
rect 1143 -723 1151 -656
rect 1217 -723 1226 -656
rect 1143 -745 1226 -723
rect 1305 -560 1397 -469
rect 1305 -642 1321 -560
rect 1378 -642 1397 -560
rect 1305 -1053 1397 -642
rect 1434 -647 1530 -328
rect 1434 -706 1447 -647
rect 1514 -706 1530 -647
rect 1434 -745 1530 -706
rect 1599 -664 1702 360
rect 1953 246 2049 263
rect 1953 193 1965 246
rect 2033 193 2049 246
rect 1953 -278 2049 193
rect 2332 -152 2420 505
rect 2331 -266 2420 -152
rect 2472 38 2560 46
rect 2472 -37 2481 38
rect 2553 -37 2560 38
rect 2472 -159 2560 -37
rect 1953 -331 1963 -278
rect 2042 -331 2049 -278
rect 1953 -333 2049 -331
rect 2332 -378 2420 -266
rect 2471 -273 2560 -159
rect 2332 -453 2338 -378
rect 2410 -453 2420 -378
rect 2332 -464 2420 -453
rect 1599 -719 1614 -664
rect 1686 -719 1702 -664
rect 1599 -745 1702 -719
rect 2076 -739 2129 -694
rect 2076 -1032 2129 -792
rect 2472 -922 2560 -273
rect 2472 -997 2481 -922
rect 2553 -997 2560 -922
rect 2472 -1009 2560 -997
rect 1305 -1111 1314 -1053
rect 1385 -1111 1397 -1053
rect 1305 -1125 1397 -1111
rect 2075 -1055 2129 -1032
rect 2075 -1109 2077 -1055
rect 2075 -1123 2129 -1109
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_0
timestamp 1746113014
transform 1 0 954 0 1 -960
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_1
timestamp 1746113014
transform 1 0 1414 0 1 -960
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  sky130_fd_sc_hd__or2_1_0
timestamp 1746113014
transform 1 0 1874 0 1 -960
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_0
timestamp 1746113014
transform 1 0 998 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_1
timestamp 1746113014
transform 1 0 1642 0 1 0
box -38 -48 682 592
<< labels >>
rlabel metal1 873 -106 873 -106 1 inA
port 1 n
rlabel metal1 869 -203 869 -203 1 inB
port 2 n
rlabel metal1 868 -312 868 -312 1 inC
port 3 n
rlabel metal1 2589 390 2589 390 1 sum
port 4 n
rlabel metal1 2633 -690 2633 -690 1 carry
port 5 n
rlabel metal1 2600 546 2600 546 1 VPWR
port 6 n
rlabel metal1 2604 -952 2604 -952 1 VGND
port 7 n
rlabel metal1 1876 -749 1876 -749 1 and1_out
rlabel metal1 1632 -1085 1632 -1085 1 and2_out
<< end >>
