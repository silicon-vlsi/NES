magic
tech sky130A
timestamp 1766122499
<< nmoslvt >>
rect -730 -110 -30 -10
rect 50 -110 750 -10
<< ndiff >>
rect -810 -30 -730 -10
rect -810 -90 -800 -30
rect -740 -90 -730 -30
rect -810 -110 -730 -90
rect -30 -20 50 -10
rect -30 -90 -10 -20
rect 30 -90 50 -20
rect -30 -110 50 -90
rect 750 -20 830 -10
rect 750 -90 770 -20
rect 810 -90 830 -20
rect 750 -110 830 -90
<< ndiffc >>
rect -800 -90 -740 -30
rect -10 -90 30 -20
rect 770 -90 810 -20
<< psubdiff >>
rect -930 150 940 170
rect -930 110 -900 150
rect 920 110 940 150
rect -930 90 940 110
rect -930 -180 -910 90
rect -870 -180 -850 90
rect -930 -190 -850 -180
rect 860 -180 880 90
rect 920 -180 940 90
rect 860 -190 940 -180
rect -930 -210 940 -190
rect -930 -250 -910 -210
rect 920 -250 940 -210
rect -930 -270 940 -250
<< psubdiffcont >>
rect -900 110 920 150
rect -910 -180 -870 90
rect 880 -180 920 90
rect -910 -250 920 -210
<< poly >>
rect -730 40 -30 60
rect -730 10 -700 40
rect -40 10 -30 40
rect -730 -10 -30 10
rect 50 40 750 60
rect 50 10 80 40
rect 740 10 750 40
rect 50 -10 750 10
rect -730 -170 -30 -110
rect 50 -170 750 -110
<< polycont >>
rect -700 10 -40 40
rect 80 10 740 40
<< locali >>
rect -920 150 930 160
rect -920 110 -900 150
rect 920 110 930 150
rect -920 100 930 110
rect -920 90 -860 100
rect -920 -180 -910 90
rect -870 -20 -860 90
rect 870 90 930 100
rect -710 40 40 50
rect -710 10 -700 40
rect -40 10 40 40
rect -710 0 40 10
rect 70 40 820 50
rect 70 10 80 40
rect 740 10 820 40
rect 70 0 820 10
rect -20 -20 40 0
rect -870 -30 -730 -20
rect -870 -90 -800 -30
rect -740 -90 -730 -30
rect -870 -100 -730 -90
rect -20 -90 -10 -20
rect 30 -90 40 -20
rect -20 -100 40 -90
rect 760 -20 820 0
rect 760 -90 770 -20
rect 810 -90 820 -20
rect 760 -100 820 -90
rect -870 -180 -860 -100
rect -920 -200 -860 -180
rect 870 -180 880 90
rect 920 -180 930 90
rect 870 -200 930 -180
rect -920 -210 930 -200
rect -920 -250 -910 -210
rect 920 -250 930 -210
rect -920 -260 930 -250
<< viali >>
rect 770 -80 810 -30
<< metal1 >>
rect 760 -30 1040 -20
rect 760 -80 770 -30
rect 810 -80 1040 -30
rect 760 -100 1040 -80
<< labels >>
rlabel psubdiffcont 30 -220 30 -220 1 gnd
port 2 n
rlabel metal1 990 -60 990 -60 1 pmosterminal
port 1 n
<< end >>
