magic
tech sky130A
timestamp 1764841088
<< pwell >>
rect 110 -235 261 958
rect 290 -235 441 958
rect 465 -235 616 958
rect 640 -235 791 958
rect 815 -235 966 958
rect 990 -235 1141 958
rect 1165 -235 1316 958
rect 1345 -235 1496 958
rect 1520 -235 1671 958
rect 1695 -235 1846 958
rect 1870 -235 2021 958
rect 2045 35 2196 958
rect 2045 -235 2195 35
rect 2220 -235 2371 958
rect 110 -1735 261 -542
rect 290 -1735 441 -542
rect 465 -1735 616 -542
rect 640 -550 645 -542
rect 1355 -550 1496 -542
rect 640 -1735 791 -550
rect 815 -1735 966 -550
rect 990 -1735 1141 -550
rect 1165 -1735 1316 -550
rect 1345 -1735 1496 -550
rect 1520 -1735 1671 -542
rect 1695 -1735 1846 -542
rect 1870 -1735 2021 -542
rect 2045 -1725 2195 -542
rect 2045 -1735 2196 -1725
rect 2220 -1735 2371 -542
<< psubdiff >>
rect -75 1305 2555 1450
rect -75 435 65 1305
rect -75 240 -50 435
rect 40 240 65 435
rect -75 -1905 65 240
rect 2415 -1905 2555 1305
rect -75 -2050 2555 -1905
<< psubdiffcont >>
rect -50 240 40 435
<< xpolycontact >>
rect 115 733 255 949
rect 115 -225 255 -9
rect 295 733 435 949
rect 295 -225 435 -9
rect 470 733 610 949
rect 470 -225 610 -9
rect 645 733 785 949
rect 645 -225 785 -9
rect 820 733 960 949
rect 820 -225 960 -9
rect 995 733 1135 949
rect 995 -225 1135 -9
rect 1170 733 1310 949
rect 1170 -225 1310 -9
rect 1350 733 1490 949
rect 1350 -225 1490 -9
rect 1525 733 1665 949
rect 1525 -225 1665 -9
rect 1700 733 1840 949
rect 1700 -225 1840 -9
rect 1875 733 2015 949
rect 1875 -225 2015 -9
rect 2050 733 2190 949
rect 2050 -225 2190 -9
rect 2225 733 2365 949
rect 2225 -225 2365 -9
rect 115 -767 255 -551
rect 115 -1725 255 -1509
rect 295 -767 435 -551
rect 295 -1725 435 -1509
rect 470 -767 610 -551
rect 470 -1725 610 -1509
rect 645 -767 785 -551
rect 645 -1725 785 -1509
rect 820 -767 960 -551
rect 820 -1725 960 -1509
rect 995 -767 1135 -551
rect 995 -1725 1135 -1509
rect 1170 -767 1310 -551
rect 1170 -1725 1310 -1509
rect 1350 -767 1490 -551
rect 1350 -1725 1490 -1509
rect 1525 -767 1665 -551
rect 1525 -1725 1665 -1509
rect 1700 -767 1840 -551
rect 1700 -1725 1840 -1509
rect 1875 -767 2015 -551
rect 1875 -1725 2015 -1509
rect 2050 -767 2190 -551
rect 2050 -1725 2190 -1509
rect 2225 -767 2365 -551
rect 2225 -1725 2365 -1509
<< ppolyres >>
rect 115 -9 255 733
rect 295 -9 435 733
rect 470 -9 610 733
rect 645 -9 785 733
rect 820 -9 960 733
rect 995 -9 1135 733
rect 1170 -9 1310 733
rect 1350 -9 1490 733
rect 1525 -9 1665 733
rect 1700 -9 1840 733
rect 1875 -9 2015 733
rect 2050 -9 2190 733
rect 2225 -9 2365 733
rect 115 -1509 255 -767
rect 295 -1509 435 -767
rect 470 -1509 610 -767
rect 645 -1509 785 -767
rect 820 -1509 960 -767
rect 995 -1509 1135 -767
rect 1170 -1509 1310 -767
rect 1350 -1509 1490 -767
rect 1525 -1509 1665 -767
rect 1700 -1509 1840 -767
rect 1875 -1509 2015 -767
rect 2050 -1509 2190 -767
rect 2225 -1509 2365 -767
<< locali >>
rect -65 1440 2543 1442
rect -65 1312 2545 1440
rect -65 949 55 1312
rect 295 1270 437 1280
rect 295 1155 305 1270
rect 425 1155 437 1270
rect 295 1145 437 1155
rect 294 949 437 1145
rect 820 1100 960 1110
rect 820 995 830 1100
rect 950 995 960 1100
rect -65 736 115 949
rect -65 435 55 736
rect 255 736 257 949
rect 294 733 295 949
rect 435 733 437 949
rect 470 949 785 950
rect 610 735 645 949
rect 820 949 960 995
rect 1525 1100 1665 1109
rect 1525 995 1535 1100
rect 1655 995 1665 1100
rect 995 949 1310 950
rect 1525 949 1665 995
rect 2425 951 2545 1312
rect 1875 949 2190 950
rect 2227 949 2545 951
rect 1135 735 1170 949
rect 2015 735 2050 949
rect 2365 733 2545 949
rect -65 240 -50 435
rect 40 240 55 435
rect -65 -11 55 240
rect 2425 -9 2545 733
rect -65 -222 115 -11
rect -65 -550 55 -222
rect 435 -225 470 -10
rect 645 -260 785 -225
rect 995 -260 1135 -225
rect 645 -380 1135 -260
rect 1170 -230 1310 -225
rect 1350 -230 1490 -225
rect 1170 -380 1490 -230
rect 1840 -225 1875 -10
rect 2365 -225 2545 -9
rect 820 -415 960 -400
rect 820 -505 835 -415
rect 945 -505 960 -415
rect -65 -551 255 -550
rect -65 -765 115 -551
rect -65 -1514 55 -765
rect 295 -551 785 -550
rect 435 -765 470 -551
rect 610 -765 645 -551
rect 820 -551 960 -505
rect 995 -551 1310 -550
rect 1525 -551 1665 -225
rect 1714 -407 2382 -399
rect 1714 -516 1723 -407
rect 1883 -414 2382 -407
rect 1883 -512 2240 -414
rect 2365 -512 2382 -414
rect 1883 -516 2382 -512
rect 1714 -526 2382 -516
rect 2425 -550 2545 -225
rect 1875 -551 2190 -550
rect 2227 -551 2545 -550
rect 1135 -765 1170 -551
rect 2015 -765 2050 -551
rect 2365 -767 2545 -551
rect 2227 -768 2545 -767
rect -65 -1722 115 -1514
rect -65 -1915 55 -1722
rect 255 -1722 257 -1514
rect 435 -1725 470 -1510
rect 1310 -1725 1350 -1510
rect 1840 -1725 1875 -1510
rect 2425 -1510 2545 -768
rect 2365 -1725 2545 -1510
rect 295 -1750 435 -1725
rect 295 -1870 305 -1750
rect 425 -1870 435 -1750
rect 295 -1880 435 -1870
rect 645 -1750 785 -1725
rect 995 -1750 1135 -1725
rect 2226 -1728 2545 -1725
rect 645 -1885 1135 -1750
rect 2425 -1915 2545 -1728
rect -65 -2040 2545 -1915
<< viali >>
rect 305 1155 425 1270
rect 830 995 950 1100
rect 1535 995 1655 1100
rect 1360 745 1480 940
rect 1710 745 1830 940
rect 830 -205 945 -30
rect 1537 -204 1656 -23
rect 2060 -215 2180 -20
rect 835 -505 945 -415
rect 1723 -516 1883 -407
rect 2240 -512 2365 -414
rect 1359 -758 1483 -560
rect 1707 -758 1831 -560
rect 835 -1710 945 -1525
rect 1540 -1710 1650 -1525
rect 2060 -1715 2180 -1520
rect 305 -1870 425 -1750
<< metal1 >>
rect -105 1270 437 1280
rect -105 1155 305 1270
rect 425 1155 437 1270
rect -105 1145 437 1155
rect -105 1109 -81 1110
rect -105 1100 1665 1109
rect -105 995 830 1100
rect 950 995 1535 1100
rect 1655 995 1665 1100
rect -105 984 1665 995
rect 1350 940 1840 950
rect 1350 745 1360 940
rect 1480 745 1710 940
rect 1830 745 1840 940
rect 1350 735 1840 745
rect 820 -23 1665 -10
rect 820 -30 1537 -23
rect 820 -205 830 -30
rect 945 -204 1537 -30
rect 1656 -204 1665 -23
rect 945 -205 1665 -204
rect 820 -225 1665 -205
rect 2050 -20 2190 -10
rect 2050 -215 2060 -20
rect 2180 -215 2190 -20
rect 727 -400 1896 -399
rect -88 -407 1896 -400
rect -88 -415 1723 -407
rect -88 -505 835 -415
rect 945 -505 1723 -415
rect -88 -516 1723 -505
rect 1883 -516 1896 -407
rect -88 -525 1896 -516
rect 1350 -560 1840 -551
rect 1350 -758 1359 -560
rect 1483 -758 1707 -560
rect 1831 -758 1840 -560
rect 1350 -766 1840 -758
rect 820 -1525 1665 -1510
rect 820 -1710 835 -1525
rect 945 -1710 1540 -1525
rect 1650 -1710 1665 -1525
rect 820 -1725 1665 -1710
rect 2050 -1520 2190 -215
rect 2223 -414 2597 -398
rect 2223 -512 2240 -414
rect 2365 -512 2597 -414
rect 2223 -525 2597 -512
rect 2050 -1715 2060 -1520
rect 2180 -1715 2190 -1520
rect 2050 -1725 2190 -1715
rect -100 -1750 435 -1740
rect -100 -1870 305 -1750
rect 425 -1870 435 -1750
rect -100 -1885 435 -1870
<< end >>
