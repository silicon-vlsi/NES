magic
tech sky130A
timestamp 1767953252
<< nwell >>
rect -20 135 165 315
<< nmos >>
rect 45 51 60 93
rect 90 51 105 93
<< pmos >>
rect 45 160 60 219
rect 90 160 105 219
<< ndiff >>
rect 18 79 45 93
rect 18 62 22 79
rect 39 62 45 79
rect 18 51 45 62
rect 60 79 90 93
rect 60 62 66 79
rect 84 62 90 79
rect 60 51 90 62
rect 105 79 133 93
rect 105 62 111 79
rect 129 62 133 79
rect 105 51 133 62
<< pdiff >>
rect 18 211 45 219
rect 18 194 22 211
rect 39 194 45 211
rect 18 160 45 194
rect 60 211 90 219
rect 60 194 66 211
rect 84 194 90 211
rect 60 160 90 194
rect 105 211 135 219
rect 105 194 111 211
rect 129 194 135 211
rect 105 160 135 194
<< ndiffc >>
rect 22 62 39 79
rect 66 62 84 79
rect 111 62 129 79
<< pdiffc >>
rect 22 194 39 211
rect 66 194 84 211
rect 111 194 129 211
<< psubdiff >>
rect 0 7 144 24
rect 0 -10 15 7
rect 32 -10 65 7
rect 82 -10 111 7
rect 129 -10 144 7
rect 0 -24 144 -10
<< nsubdiff >>
rect 0 278 146 295
rect 0 261 15 278
rect 32 261 65 278
rect 82 261 111 278
rect 129 261 146 278
rect 0 246 146 261
<< psubdiffcont >>
rect 15 -10 32 7
rect 65 -10 82 7
rect 111 -10 129 7
<< nsubdiffcont >>
rect 15 261 32 278
rect 65 261 82 278
rect 111 261 129 278
<< poly >>
rect 45 219 60 232
rect 90 219 105 232
rect 45 143 60 160
rect 15 135 60 143
rect 15 118 20 135
rect 37 118 60 135
rect 15 110 60 118
rect 45 93 60 110
rect 90 143 105 160
rect 90 135 135 143
rect 90 118 110 135
rect 127 118 135 135
rect 90 110 135 118
rect 90 93 105 110
rect 45 38 60 51
rect 90 38 105 51
<< polycont >>
rect 20 118 37 135
rect 110 118 127 135
<< locali >>
rect 0 278 146 295
rect 0 261 15 278
rect 32 261 65 278
rect 82 261 111 278
rect 129 261 146 278
rect 0 246 146 261
rect 18 211 43 246
rect 63 219 88 220
rect 18 194 22 211
rect 39 194 43 211
rect 18 160 43 194
rect 62 211 88 219
rect 62 194 66 211
rect 84 194 88 211
rect 62 160 88 194
rect 107 211 135 219
rect 107 194 111 211
rect 129 194 135 211
rect 107 160 135 194
rect 15 135 45 143
rect 15 118 20 135
rect 37 118 45 135
rect 15 110 45 118
rect 105 135 135 143
rect 105 118 110 135
rect 127 118 135 135
rect 105 110 135 118
rect 18 79 43 93
rect 18 62 22 79
rect 39 62 43 79
rect 18 24 43 62
rect 62 79 88 93
rect 62 62 66 79
rect 84 62 88 79
rect 62 51 88 62
rect 107 79 133 93
rect 107 62 111 79
rect 129 62 133 79
rect 107 51 133 62
rect 63 50 88 51
rect 108 24 133 51
rect 0 7 144 24
rect 0 -10 15 7
rect 32 -10 65 7
rect 82 -10 111 7
rect 129 -10 144 7
rect 0 -25 144 -10
<< viali >>
rect 15 261 32 278
rect 65 261 82 278
rect 111 261 129 278
rect 111 194 129 211
rect 20 118 37 135
rect 110 118 127 135
rect 66 62 84 79
rect 15 -10 32 7
rect 65 -10 82 7
rect 111 -10 129 7
<< metal1 >>
rect 0 278 146 295
rect 0 261 15 278
rect 32 261 65 278
rect 82 261 111 278
rect 129 261 146 278
rect 0 246 146 261
rect 62 211 136 215
rect 62 194 111 211
rect 129 194 136 211
rect 62 190 136 194
rect 15 142 45 143
rect 15 135 46 142
rect 15 118 20 135
rect 37 118 46 135
rect 15 111 46 118
rect 15 110 45 111
rect 62 79 88 190
rect 105 135 135 143
rect 105 118 110 135
rect 127 118 135 135
rect 105 110 135 118
rect 62 62 66 79
rect 84 65 88 79
rect 84 62 87 65
rect 62 52 87 62
rect 0 7 144 24
rect 0 -10 15 7
rect 32 -10 65 7
rect 82 -10 111 7
rect 129 -10 144 7
rect 0 -25 144 -10
<< labels >>
rlabel nwell 9 256 137 287 1 vdd
port 1 n
rlabel metal1 11 -16 139 15 1 gnd
port 2 n
rlabel metal1 109 114 131 132 1 b
port 3 n
rlabel metal1 20 114 42 132 1 a
port 4 n
rlabel metal1 65 110 87 128 1 out
port 5 n
<< end >>
