magic
tech sky130A
timestamp 1767782451
<< fence >>
rect 0 0 245 270
<< nwell >>
rect -20 135 265 315
<< nmos >>
rect 45 51 60 93
rect 90 51 105 93
rect 140 51 155 93
rect 185 51 200 93
<< pmos >>
rect 45 160 60 219
rect 90 160 105 219
rect 140 160 155 219
rect 185 160 200 219
<< ndiff >>
rect 18 79 45 93
rect 18 62 22 79
rect 39 62 45 79
rect 18 51 45 62
rect 60 79 90 93
rect 60 62 66 79
rect 84 62 90 79
rect 60 51 90 62
rect 105 79 140 93
rect 105 62 111 79
rect 134 62 140 79
rect 105 51 140 62
rect 155 79 185 93
rect 155 62 161 79
rect 179 62 185 79
rect 155 51 185 62
rect 200 79 227 93
rect 200 62 206 79
rect 223 62 227 79
rect 200 51 227 62
<< pdiff >>
rect 18 211 45 219
rect 18 194 22 211
rect 39 194 45 211
rect 18 160 45 194
rect 60 211 90 219
rect 60 194 66 211
rect 84 194 90 211
rect 60 160 90 194
rect 105 211 140 219
rect 105 194 111 211
rect 134 194 140 211
rect 105 160 140 194
rect 155 211 185 219
rect 155 194 161 211
rect 179 194 185 211
rect 155 160 185 194
rect 200 211 227 219
rect 200 194 206 211
rect 223 194 227 211
rect 200 160 227 194
<< ndiffc >>
rect 22 62 39 79
rect 66 62 84 79
rect 111 62 134 79
rect 161 62 179 79
rect 206 62 223 79
<< pdiffc >>
rect 22 194 39 211
rect 66 194 84 211
rect 111 194 134 211
rect 161 194 179 211
rect 206 194 223 211
<< psubdiff >>
rect 0 7 245 24
rect 0 -10 15 7
rect 32 -10 66 7
rect 84 -10 112 7
rect 132 -10 161 7
rect 179 -10 213 7
rect 230 -10 245 7
rect 0 -24 245 -10
<< nsubdiff >>
rect 0 278 245 294
rect 0 261 15 278
rect 32 261 66 278
rect 84 261 110 278
rect 130 261 161 278
rect 179 261 213 278
rect 230 261 245 278
rect 0 246 245 261
<< psubdiffcont >>
rect 15 -10 32 7
rect 66 -10 84 7
rect 112 -10 132 7
rect 161 -10 179 7
rect 213 -10 230 7
<< nsubdiffcont >>
rect 15 261 32 278
rect 66 261 84 278
rect 110 261 130 278
rect 161 261 179 278
rect 213 261 230 278
<< poly >>
rect 45 219 60 232
rect 90 219 105 232
rect 140 219 155 232
rect 185 219 200 232
rect 45 143 60 160
rect 15 135 60 143
rect 15 118 20 135
rect 37 118 60 135
rect 15 110 60 118
rect 45 93 60 110
rect 90 143 105 160
rect 140 143 155 160
rect 90 135 155 143
rect 90 118 113 135
rect 132 118 155 135
rect 90 110 155 118
rect 90 93 105 110
rect 140 93 155 110
rect 185 143 200 160
rect 185 135 230 143
rect 185 118 208 135
rect 225 118 230 135
rect 185 110 230 118
rect 185 93 200 110
rect 45 38 60 51
rect 90 38 105 51
rect 140 38 155 51
rect 185 38 200 51
<< polycont >>
rect 20 118 37 135
rect 113 118 132 135
rect 208 118 225 135
<< locali >>
rect 0 278 245 295
rect 0 261 15 278
rect 32 261 66 278
rect 84 261 110 278
rect 130 261 161 278
rect 179 261 213 278
rect 230 261 245 278
rect 0 245 245 261
rect 18 211 43 245
rect 18 194 22 211
rect 39 194 43 211
rect 18 160 43 194
rect 62 211 88 219
rect 62 194 66 211
rect 84 194 88 211
rect 15 135 45 143
rect 15 118 20 135
rect 37 118 45 135
rect 15 110 45 118
rect 18 79 43 93
rect 18 62 22 79
rect 39 62 43 79
rect 18 24 43 62
rect 62 79 88 194
rect 107 211 138 245
rect 107 194 111 211
rect 134 194 138 211
rect 107 160 138 194
rect 157 211 183 219
rect 157 194 161 211
rect 179 194 183 211
rect 105 135 140 143
rect 105 118 113 135
rect 132 118 140 135
rect 105 110 140 118
rect 62 62 66 79
rect 84 62 88 79
rect 62 51 88 62
rect 107 79 138 93
rect 107 62 111 79
rect 134 62 138 79
rect 107 24 138 62
rect 157 79 183 194
rect 202 211 227 245
rect 202 194 206 211
rect 223 194 227 211
rect 202 160 227 194
rect 200 135 230 143
rect 200 118 208 135
rect 225 118 230 135
rect 200 110 230 118
rect 157 62 161 79
rect 179 62 183 79
rect 157 51 183 62
rect 202 79 227 93
rect 202 62 206 79
rect 223 62 227 79
rect 202 24 227 62
rect 0 7 245 24
rect 0 -10 15 7
rect 32 -10 66 7
rect 84 -10 112 7
rect 132 -10 161 7
rect 179 -10 213 7
rect 230 -10 245 7
rect 0 -25 245 -10
<< viali >>
rect 15 261 32 278
rect 66 261 84 278
rect 110 261 130 278
rect 161 261 179 278
rect 213 261 230 278
rect 66 194 84 211
rect 20 118 37 135
rect 161 194 179 211
rect 113 118 132 135
rect 208 118 225 135
rect 15 -10 32 7
rect 66 -10 84 7
rect 112 -10 132 7
rect 161 -10 179 7
rect 213 -10 230 7
<< metal1 >>
rect 0 278 245 295
rect 0 261 15 278
rect 32 261 66 278
rect 84 261 110 278
rect 130 261 161 278
rect 179 261 213 278
rect 230 261 245 278
rect 0 245 245 261
rect 60 211 186 217
rect 60 194 66 211
rect 84 194 161 211
rect 179 194 186 211
rect 60 185 186 194
rect 15 142 45 143
rect 105 142 140 143
rect 200 142 230 143
rect 15 135 231 142
rect 15 118 20 135
rect 37 118 113 135
rect 132 118 208 135
rect 225 118 231 135
rect 15 111 231 118
rect 15 110 45 111
rect 105 110 140 111
rect 200 110 230 111
rect 0 7 245 24
rect 0 -10 15 7
rect 32 -10 66 7
rect 84 -10 112 7
rect 132 -10 161 7
rect 179 -10 213 7
rect 230 -10 245 7
rect 0 -25 245 -10
<< labels >>
rlabel nwell 10 256 235 284 1 vdd
port 1 n
rlabel metal1 11 -16 236 12 1 gnd
port 2 n
rlabel metal1 204 112 228 133 1 in
port 3 n
rlabel locali 163 97 182 104 1 out
port 4 n
<< end >>
