magic
tech sky130A
timestamp 1766123683
<< nmoslvt >>
rect -60 200 40 700
rect 140 200 240 700
rect 340 200 440 700
rect 540 200 640 700
rect 740 200 840 700
rect 940 200 1040 700
rect 1140 200 1240 700
rect 1340 200 1440 700
rect 1540 200 1640 700
rect 1740 200 1840 700
rect 1940 200 2040 700
rect 2140 200 2240 700
rect 2340 200 2440 700
rect 2540 200 2640 700
rect -60 -770 40 -270
rect 140 -770 240 -270
rect 340 -770 440 -270
rect 540 -770 640 -270
rect 740 -770 840 -270
rect 940 -770 1040 -270
rect 1140 -770 1240 -270
rect 1340 -770 1440 -270
rect 1540 -770 1640 -270
rect 1740 -770 1840 -270
rect 1940 -770 2040 -270
rect 2140 -770 2240 -270
rect 2340 -770 2440 -270
rect 2540 -770 2640 -270
<< ndiff >>
rect -160 690 -60 700
rect -160 470 -140 690
rect -80 470 -60 690
rect -160 200 -60 470
rect 40 440 140 700
rect 40 220 60 440
rect 120 220 140 440
rect 40 200 140 220
rect 240 690 340 700
rect 240 470 260 690
rect 320 470 340 690
rect 240 200 340 470
rect 440 440 540 700
rect 440 220 460 440
rect 520 220 540 440
rect 440 200 540 220
rect 640 690 740 700
rect 640 490 660 690
rect 720 490 740 690
rect 640 200 740 490
rect 840 690 940 700
rect 840 490 860 690
rect 920 490 940 690
rect 840 200 940 490
rect 1040 430 1140 700
rect 1040 230 1060 430
rect 1120 230 1140 430
rect 1040 200 1140 230
rect 1240 690 1340 700
rect 1240 490 1260 690
rect 1320 490 1340 690
rect 1240 200 1340 490
rect 1440 430 1540 700
rect 1440 230 1460 430
rect 1520 230 1540 430
rect 1440 200 1540 230
rect 1640 690 1740 700
rect 1640 490 1660 690
rect 1720 490 1740 690
rect 1640 200 1740 490
rect 1840 690 1940 700
rect 1840 480 1860 690
rect 1920 480 1940 690
rect 1840 200 1940 480
rect 2040 440 2140 700
rect 2040 210 2060 440
rect 2120 210 2140 440
rect 2040 200 2140 210
rect 2240 690 2340 700
rect 2240 460 2260 690
rect 2320 460 2340 690
rect 2240 200 2340 460
rect 2440 440 2540 700
rect 2440 210 2460 440
rect 2520 210 2540 440
rect 2440 200 2540 210
rect 2640 690 2740 700
rect 2640 470 2660 690
rect 2720 470 2740 690
rect 2640 200 2740 470
rect -160 -520 -60 -270
rect -160 -760 -140 -520
rect -80 -760 -60 -520
rect -160 -770 -60 -760
rect 40 -530 140 -270
rect 40 -750 60 -530
rect 120 -750 140 -530
rect 40 -770 140 -750
rect 240 -280 340 -270
rect 240 -500 260 -280
rect 320 -500 340 -280
rect 240 -770 340 -500
rect 440 -530 540 -270
rect 440 -750 460 -530
rect 520 -750 540 -530
rect 440 -770 540 -750
rect 640 -520 740 -270
rect 640 -760 660 -520
rect 720 -760 740 -520
rect 640 -770 740 -760
rect 840 -490 940 -270
rect 840 -760 860 -490
rect 920 -760 940 -490
rect 840 -770 940 -760
rect 1040 -280 1140 -270
rect 1040 -540 1060 -280
rect 1120 -540 1140 -280
rect 1040 -770 1140 -540
rect 1240 -490 1340 -270
rect 1240 -760 1260 -490
rect 1320 -760 1340 -490
rect 1240 -770 1340 -760
rect 1440 -280 1540 -270
rect 1440 -540 1460 -280
rect 1520 -540 1540 -280
rect 1440 -770 1540 -540
rect 1640 -490 1740 -270
rect 1640 -760 1660 -490
rect 1720 -760 1740 -490
rect 1640 -770 1740 -760
rect 1840 -530 1940 -270
rect 1840 -760 1860 -530
rect 1920 -760 1940 -530
rect 1840 -770 1940 -760
rect 2040 -530 2140 -270
rect 2040 -760 2060 -530
rect 2120 -760 2140 -530
rect 2040 -770 2140 -760
rect 2240 -280 2340 -270
rect 2240 -500 2260 -280
rect 2320 -500 2340 -280
rect 2240 -770 2340 -500
rect 2440 -530 2540 -270
rect 2440 -750 2460 -530
rect 2520 -750 2540 -530
rect 2440 -770 2540 -750
rect 2640 -520 2740 -270
rect 2640 -760 2660 -520
rect 2720 -760 2740 -520
rect 2640 -770 2740 -760
<< ndiffc >>
rect -140 470 -80 690
rect 60 220 120 440
rect 260 470 320 690
rect 460 220 520 440
rect 660 490 720 690
rect 860 490 920 690
rect 1060 230 1120 430
rect 1260 490 1320 690
rect 1460 230 1520 430
rect 1660 490 1720 690
rect 1860 480 1920 690
rect 2060 210 2120 440
rect 2260 460 2320 690
rect 2460 210 2520 440
rect 2660 470 2720 690
rect -140 -760 -80 -520
rect 60 -750 120 -530
rect 260 -500 320 -280
rect 460 -750 520 -530
rect 660 -760 720 -520
rect 860 -760 920 -490
rect 1060 -540 1120 -280
rect 1260 -760 1320 -490
rect 1460 -540 1520 -280
rect 1660 -760 1720 -490
rect 1860 -760 1920 -530
rect 2060 -760 2120 -530
rect 2260 -500 2320 -280
rect 2460 -750 2520 -530
rect 2660 -760 2720 -520
<< psubdiff >>
rect -300 1150 3200 1170
rect -300 690 -280 1150
rect -210 1080 -140 1150
rect 640 1080 660 1150
rect -210 1070 660 1080
rect 1920 1070 1950 1150
rect 2720 1070 3200 1150
rect -210 1050 3200 1070
rect -210 690 -190 1050
rect 3090 780 3200 1050
rect -300 620 -190 690
rect -300 160 -280 620
rect -210 160 -190 620
rect 3090 310 3110 780
rect 3180 310 3200 780
rect -300 40 -190 160
rect -300 -420 -280 40
rect -210 -420 -190 40
rect 3090 -200 3200 310
rect -300 -760 -190 -420
rect -300 -1220 -280 -760
rect -210 -1150 -190 -760
rect 3090 -670 3110 -200
rect 3180 -670 3200 -200
rect 3090 -1150 3200 -670
rect -210 -1170 3200 -1150
rect -210 -1220 -180 -1170
rect -300 -1250 -180 -1220
rect 850 -1250 970 -1170
rect 2000 -1250 2090 -1170
rect 3140 -1250 3200 -1170
rect -300 -1270 3200 -1250
<< psubdiffcont >>
rect -280 690 -210 1150
rect -140 1080 640 1150
rect 660 1070 1920 1150
rect 1950 1070 2720 1150
rect -280 160 -210 620
rect 3110 310 3180 780
rect -280 -420 -210 40
rect -280 -1220 -210 -760
rect 3110 -670 3180 -200
rect -180 -1250 850 -1170
rect 970 -1250 2000 -1170
rect 2090 -1250 3140 -1170
<< poly >>
rect 140 890 240 900
rect 140 800 150 890
rect 220 800 240 890
rect -60 770 40 790
rect -60 720 -50 770
rect 30 720 40 770
rect -60 700 40 720
rect 140 700 240 800
rect 340 890 440 900
rect 340 800 360 890
rect 430 800 440 890
rect 340 700 440 800
rect 2140 890 2240 900
rect 2140 800 2150 890
rect 2220 800 2240 890
rect 540 750 640 770
rect 540 720 560 750
rect 630 720 640 750
rect 540 700 640 720
rect 740 750 840 770
rect 740 720 750 750
rect 820 720 840 750
rect 740 700 840 720
rect 940 760 1040 770
rect 940 720 960 760
rect 1020 720 1040 760
rect 940 700 1040 720
rect 1140 760 1240 770
rect 1140 720 1160 760
rect 1220 720 1240 760
rect 1140 700 1240 720
rect 1340 760 1440 770
rect 1340 720 1360 760
rect 1420 720 1440 760
rect 1340 700 1440 720
rect 1540 760 1640 770
rect 1540 720 1560 760
rect 1620 720 1640 760
rect 1540 700 1640 720
rect 1740 750 1840 770
rect 1740 720 1760 750
rect 1830 720 1840 750
rect 1740 700 1840 720
rect 1940 750 2040 770
rect 1940 720 1950 750
rect 2020 720 2040 750
rect 1940 700 2040 720
rect 2140 700 2240 800
rect 2340 890 2440 900
rect 2340 800 2350 890
rect 2430 800 2440 890
rect 2340 700 2440 800
rect 2540 750 2640 770
rect 2540 720 2560 750
rect 2630 720 2640 750
rect 2540 700 2640 720
rect -60 150 40 200
rect 140 150 240 200
rect 340 150 440 200
rect 540 160 640 200
rect 740 160 840 200
rect 940 150 1040 200
rect 1140 150 1240 200
rect 1340 150 1440 200
rect 1540 150 1640 200
rect 1740 150 1840 200
rect 1940 150 2040 200
rect 2140 150 2240 200
rect 2340 150 2440 200
rect 2540 160 2640 200
rect -60 -270 40 -220
rect 140 -270 240 -220
rect 340 -270 440 -220
rect 540 -270 640 -220
rect 740 -270 840 -220
rect 940 -270 1040 -200
rect 1140 -270 1240 -200
rect 1340 -270 1440 -200
rect 1540 -270 1640 -200
rect 1740 -270 1840 -200
rect 1940 -270 2040 -200
rect 2140 -270 2240 -220
rect 2340 -270 2440 -220
rect 2540 -270 2640 -220
rect -60 -790 40 -770
rect -60 -840 -50 -790
rect 20 -840 40 -790
rect -60 -850 40 -840
rect 140 -790 240 -770
rect 140 -830 160 -790
rect 230 -830 240 -790
rect 140 -850 240 -830
rect 340 -790 440 -770
rect 340 -830 350 -790
rect 420 -830 440 -790
rect 340 -850 440 -830
rect 540 -790 640 -770
rect 540 -830 560 -790
rect 630 -830 640 -790
rect 540 -850 640 -830
rect 740 -790 840 -770
rect 740 -830 750 -790
rect 820 -830 840 -790
rect 740 -850 840 -830
rect 940 -870 1040 -770
rect 940 -960 960 -870
rect 1030 -960 1040 -870
rect 940 -970 1040 -960
rect 1140 -870 1240 -770
rect 1140 -960 1150 -870
rect 1220 -960 1240 -870
rect 1140 -970 1240 -960
rect 1340 -870 1440 -770
rect 1340 -960 1360 -870
rect 1430 -960 1440 -870
rect 1340 -970 1440 -960
rect 1540 -870 1640 -770
rect 1740 -790 1840 -770
rect 1740 -830 1760 -790
rect 1830 -830 1840 -790
rect 1740 -850 1840 -830
rect 1940 -790 2040 -770
rect 1940 -830 1950 -790
rect 2020 -830 2040 -790
rect 1940 -850 2040 -830
rect 2140 -790 2240 -770
rect 2140 -830 2160 -790
rect 2230 -830 2240 -790
rect 2140 -850 2240 -830
rect 2340 -790 2440 -770
rect 2340 -830 2350 -790
rect 2420 -830 2440 -790
rect 2340 -850 2440 -830
rect 2540 -790 2640 -770
rect 2540 -830 2560 -790
rect 2630 -830 2640 -790
rect 2540 -850 2640 -830
rect 1540 -960 1550 -870
rect 1620 -960 1640 -870
rect 1540 -970 1640 -960
<< polycont >>
rect 150 800 220 890
rect -50 720 30 770
rect 360 800 430 890
rect 2150 800 2220 890
rect 560 720 630 750
rect 750 720 820 750
rect 960 720 1020 760
rect 1160 720 1220 760
rect 1360 720 1420 760
rect 1560 720 1620 760
rect 1760 720 1830 750
rect 1950 720 2020 750
rect 2350 800 2430 890
rect 2560 720 2630 750
rect -50 -840 20 -790
rect 160 -830 230 -790
rect 350 -830 420 -790
rect 560 -830 630 -790
rect 750 -830 820 -790
rect 960 -960 1030 -870
rect 1150 -960 1220 -870
rect 1360 -960 1430 -870
rect 1760 -830 1830 -790
rect 1950 -830 2020 -790
rect 2160 -830 2230 -790
rect 2350 -830 2420 -790
rect 2560 -830 2630 -790
rect 1550 -960 1620 -870
<< locali >>
rect 2650 1160 2730 1170
rect -290 1150 3190 1160
rect -290 690 -280 1150
rect -210 1080 -140 1150
rect 640 1080 660 1150
rect -210 1070 660 1080
rect 1920 1070 1950 1150
rect 2720 1070 3190 1150
rect -210 1060 3190 1070
rect -210 690 -200 1060
rect -290 620 -200 690
rect -290 160 -280 620
rect -210 160 -200 620
rect -150 780 -70 1060
rect 250 1010 330 1020
rect 250 930 260 1010
rect 320 930 330 1010
rect 140 890 230 900
rect 140 800 150 890
rect 220 800 230 890
rect 140 790 230 800
rect -150 770 40 780
rect -150 720 -50 770
rect 30 720 40 770
rect -150 710 40 720
rect -150 690 -70 710
rect -150 470 -140 690
rect -80 470 -70 690
rect -150 450 -70 470
rect 250 690 330 930
rect 350 890 440 900
rect 350 800 360 890
rect 430 800 440 890
rect 350 790 440 800
rect 650 760 730 1060
rect 850 890 930 900
rect 850 800 860 890
rect 920 800 930 890
rect 850 770 930 800
rect 1250 890 1330 900
rect 1250 800 1260 890
rect 1320 800 1330 890
rect 1250 770 1330 800
rect 1650 890 1730 900
rect 1650 800 1660 890
rect 1720 800 1730 890
rect 1650 770 1730 800
rect 850 760 1730 770
rect 1850 760 1930 1060
rect 2250 1010 2330 1020
rect 2250 930 2260 1010
rect 2320 930 2330 1010
rect 2140 890 2230 900
rect 2140 800 2150 890
rect 2220 800 2230 890
rect 2140 790 2230 800
rect 550 750 830 760
rect 550 720 560 750
rect 630 720 750 750
rect 820 720 830 750
rect 550 710 830 720
rect 850 720 960 760
rect 1020 720 1160 760
rect 1220 720 1360 760
rect 1420 720 1560 760
rect 1620 720 1730 760
rect 850 710 1730 720
rect 1750 750 2030 760
rect 1750 720 1760 750
rect 1830 720 1950 750
rect 2020 720 2030 750
rect 1750 710 2030 720
rect 250 470 260 690
rect 320 470 330 690
rect 650 690 730 710
rect 650 490 660 690
rect 720 490 730 690
rect 650 470 730 490
rect 850 690 930 710
rect 850 490 860 690
rect 920 490 930 690
rect 850 470 930 490
rect 1250 690 1330 710
rect 1250 490 1260 690
rect 1320 490 1330 690
rect 1250 470 1330 490
rect 1650 690 1730 710
rect 1650 490 1660 690
rect 1720 490 1730 690
rect 1650 470 1730 490
rect 1850 690 1930 710
rect 1850 480 1860 690
rect 1920 480 1930 690
rect 1850 470 1930 480
rect 2250 690 2330 930
rect 2350 890 2440 900
rect 2430 800 2440 890
rect 2350 790 2440 800
rect 2650 760 2730 1060
rect 2550 750 2730 760
rect 2550 720 2560 750
rect 2630 720 2730 750
rect 2550 710 2730 720
rect 250 450 330 470
rect 2250 460 2260 690
rect 2320 460 2330 690
rect 2650 690 2730 710
rect 2650 470 2660 690
rect 2720 470 2730 690
rect 2650 460 2730 470
rect 2780 1010 2900 1020
rect 2780 930 2790 1010
rect 2890 930 2900 1010
rect 2250 450 2330 460
rect -290 40 -200 160
rect -290 -420 -280 40
rect -210 -420 -200 40
rect 50 440 130 450
rect 50 220 60 440
rect 120 220 130 440
rect 50 -80 130 220
rect 450 440 530 450
rect 450 220 460 440
rect 520 220 530 440
rect 50 -170 60 -80
rect 120 -170 130 -80
rect 50 -180 130 -170
rect 250 70 330 80
rect 250 -20 260 70
rect 320 -20 330 70
rect -290 -760 -200 -420
rect 250 -280 330 -20
rect 450 -80 530 220
rect 1050 430 1130 450
rect 1050 230 1060 430
rect 1120 230 1130 430
rect 1050 70 1130 230
rect 1050 -20 1060 70
rect 1120 -20 1130 70
rect 1050 -30 1130 -20
rect 1450 430 1530 450
rect 1450 230 1460 430
rect 1520 230 1530 430
rect 1450 70 1530 230
rect 1450 -20 1460 70
rect 1520 -20 1530 70
rect 1450 -30 1530 -20
rect 2050 440 2130 450
rect 2050 210 2060 440
rect 2120 210 2130 440
rect 450 -170 460 -80
rect 520 -170 530 -80
rect 450 -180 530 -170
rect 1050 -80 1130 -70
rect 1050 -170 1060 -80
rect 1120 -170 1130 -80
rect 250 -500 260 -280
rect 320 -500 330 -280
rect 1050 -280 1130 -170
rect 250 -510 330 -500
rect 850 -490 930 -480
rect -290 -1220 -280 -760
rect -210 -1160 -200 -760
rect -150 -520 -70 -510
rect -150 -760 -140 -520
rect -80 -760 -70 -520
rect -150 -780 -70 -760
rect 50 -530 130 -510
rect 50 -750 60 -530
rect 120 -750 130 -530
rect -150 -790 30 -780
rect -150 -840 -50 -790
rect 20 -840 30 -790
rect -150 -850 30 -840
rect -150 -1160 -70 -850
rect 50 -870 130 -750
rect 450 -530 530 -510
rect 450 -750 460 -530
rect 520 -750 530 -530
rect 150 -790 430 -780
rect 150 -830 160 -790
rect 230 -830 350 -790
rect 420 -830 430 -790
rect 150 -840 430 -830
rect 50 -960 60 -870
rect 120 -960 130 -870
rect 50 -970 130 -960
rect 250 -870 330 -840
rect 250 -960 260 -870
rect 320 -960 330 -870
rect 250 -970 330 -960
rect 450 -870 530 -750
rect 650 -520 730 -510
rect 650 -760 660 -520
rect 720 -760 730 -520
rect 650 -780 730 -760
rect 850 -760 860 -490
rect 920 -760 930 -490
rect 1050 -540 1060 -280
rect 1120 -540 1130 -280
rect 1450 -80 1530 -70
rect 1450 -170 1460 -80
rect 1520 -170 1530 -80
rect 1450 -280 1530 -170
rect 2050 -80 2130 210
rect 2450 440 2530 450
rect 2450 210 2460 440
rect 2520 210 2530 440
rect 2050 -170 2060 -80
rect 2120 -170 2130 -80
rect 2050 -180 2130 -170
rect 2260 70 2340 80
rect 2260 -20 2270 70
rect 2330 -20 2340 70
rect 2260 -180 2340 -20
rect 2450 -80 2530 210
rect 2450 -170 2460 -80
rect 2520 -170 2530 -80
rect 2450 -180 2530 -170
rect 1050 -550 1130 -540
rect 1250 -490 1330 -480
rect 550 -790 830 -780
rect 550 -830 560 -790
rect 630 -830 750 -790
rect 820 -830 830 -790
rect 550 -840 830 -830
rect 450 -960 460 -870
rect 520 -960 530 -870
rect 450 -970 530 -960
rect 650 -1160 730 -840
rect 850 -1030 930 -760
rect 1250 -760 1260 -490
rect 1320 -760 1330 -490
rect 1450 -540 1460 -280
rect 1520 -540 1530 -280
rect 2250 -280 2330 -180
rect 1450 -550 1530 -540
rect 1650 -490 1730 -480
rect 950 -870 1040 -860
rect 950 -960 960 -870
rect 1030 -960 1040 -870
rect 950 -970 1040 -960
rect 1140 -870 1230 -860
rect 1140 -960 1150 -870
rect 1220 -960 1230 -870
rect 1140 -970 1230 -960
rect 850 -1120 860 -1030
rect 920 -1120 930 -1030
rect 850 -1130 930 -1120
rect 1250 -1030 1330 -760
rect 1650 -760 1660 -490
rect 1720 -760 1730 -490
rect 2250 -500 2260 -280
rect 2320 -500 2330 -280
rect 2250 -510 2330 -500
rect 1350 -870 1440 -860
rect 1350 -960 1360 -870
rect 1430 -960 1440 -870
rect 1350 -970 1440 -960
rect 1540 -870 1630 -860
rect 1540 -960 1550 -870
rect 1620 -960 1630 -870
rect 1540 -970 1630 -960
rect 1250 -1120 1260 -1030
rect 1320 -1120 1330 -1030
rect 1250 -1130 1330 -1120
rect 1650 -1030 1730 -760
rect 1850 -530 1930 -510
rect 1850 -760 1860 -530
rect 1920 -760 1930 -530
rect 1850 -780 1930 -760
rect 2050 -530 2130 -510
rect 2050 -760 2060 -530
rect 2120 -760 2130 -530
rect 1750 -790 2030 -780
rect 1750 -830 1760 -790
rect 1830 -830 1950 -790
rect 2020 -830 2030 -790
rect 1750 -840 2030 -830
rect 1650 -1120 1660 -1030
rect 1720 -1120 1730 -1030
rect 1650 -1130 1730 -1120
rect 1850 -1160 1930 -840
rect 2050 -870 2130 -760
rect 2450 -530 2530 -510
rect 2450 -750 2460 -530
rect 2520 -750 2530 -530
rect 2150 -790 2430 -780
rect 2150 -830 2160 -790
rect 2230 -830 2350 -790
rect 2420 -830 2430 -790
rect 2150 -840 2430 -830
rect 2050 -960 2060 -870
rect 2120 -960 2130 -870
rect 2050 -970 2130 -960
rect 2250 -870 2330 -840
rect 2250 -960 2260 -870
rect 2320 -960 2330 -870
rect 2250 -970 2330 -960
rect 2450 -870 2530 -750
rect 2650 -520 2730 -510
rect 2650 -760 2660 -520
rect 2720 -760 2730 -520
rect 2650 -780 2730 -760
rect 2550 -790 2730 -780
rect 2550 -830 2560 -790
rect 2630 -830 2730 -790
rect 2550 -840 2730 -830
rect 2450 -960 2460 -870
rect 2520 -960 2530 -870
rect 2450 -970 2530 -960
rect 2650 -1160 2730 -840
rect 2780 -1030 2900 930
rect 2920 890 3060 900
rect 2920 800 2930 890
rect 3050 800 3060 890
rect 2920 -870 3060 800
rect 2920 -960 2930 -870
rect 3050 -960 3060 -870
rect 2920 -970 3060 -960
rect 3100 780 3190 1060
rect 3100 310 3110 780
rect 3180 310 3190 780
rect 3100 -200 3190 310
rect 3100 -670 3110 -200
rect 3180 -670 3190 -200
rect 2780 -1120 2790 -1030
rect 2890 -1120 2900 -1030
rect 2780 -1130 2900 -1120
rect 3100 -1160 3190 -670
rect -210 -1170 3190 -1160
rect -210 -1220 -180 -1170
rect -290 -1250 -180 -1220
rect 850 -1250 970 -1170
rect 2000 -1250 2090 -1170
rect 3140 -1250 3190 -1170
rect -290 -1260 3190 -1250
<< viali >>
rect 260 930 320 1010
rect 160 810 210 880
rect 370 810 420 880
rect 860 800 920 890
rect 1260 800 1320 890
rect 1660 800 1720 890
rect 2260 930 2320 1010
rect 2160 810 2210 880
rect 2360 810 2420 880
rect 2790 930 2890 1010
rect 60 -170 120 -80
rect 260 -20 320 70
rect 1060 -20 1120 70
rect 1460 -20 1520 70
rect 460 -170 520 -80
rect 1060 -170 1120 -80
rect 60 -960 120 -870
rect 260 -960 320 -870
rect 1460 -170 1520 -80
rect 2060 -170 2120 -80
rect 2270 -20 2330 70
rect 2460 -170 2520 -80
rect 460 -960 520 -870
rect 970 -950 1020 -880
rect 1160 -950 1210 -880
rect 860 -1120 920 -1030
rect 1370 -950 1420 -880
rect 1560 -950 1610 -880
rect 1260 -1120 1320 -1030
rect 1660 -1120 1720 -1030
rect 2060 -960 2120 -870
rect 2260 -960 2320 -870
rect 2460 -960 2520 -870
rect 2930 800 3050 890
rect 2930 -960 3050 -870
rect 2790 -1120 2890 -1030
<< metal1 >>
rect 130 1010 2920 1020
rect 130 930 260 1010
rect 320 930 2260 1010
rect 2320 930 2790 1010
rect 2890 930 2920 1010
rect 130 920 2920 930
rect 140 890 3266 900
rect 140 880 860 890
rect 140 810 160 880
rect 210 810 370 880
rect 420 810 860 880
rect 140 800 860 810
rect 920 800 1260 890
rect 1320 800 1660 890
rect 1720 880 2930 890
rect 1720 810 2160 880
rect 2210 810 2360 880
rect 2420 810 2930 880
rect 1720 800 2930 810
rect 3050 800 3266 890
rect 140 790 3266 800
rect 40 70 3266 80
rect 40 -20 260 70
rect 320 -20 1060 70
rect 1120 -20 1460 70
rect 1520 -20 2270 70
rect 2330 -20 3266 70
rect 40 -30 3266 -20
rect 40 -80 3266 -70
rect 40 -170 60 -80
rect 120 -170 460 -80
rect 520 -170 1060 -80
rect 1120 -170 1460 -80
rect 1520 -170 2060 -80
rect 2120 -170 2460 -80
rect 2520 -170 3266 -80
rect 40 -180 3266 -170
rect 40 -870 3080 -860
rect 40 -960 60 -870
rect 120 -960 260 -870
rect 320 -960 460 -870
rect 520 -880 2060 -870
rect 520 -950 970 -880
rect 1020 -950 1160 -880
rect 1210 -950 1370 -880
rect 1420 -950 1560 -880
rect 1610 -950 2060 -880
rect 520 -960 2060 -950
rect 2120 -960 2260 -870
rect 2320 -960 2460 -870
rect 2520 -960 2930 -870
rect 3050 -960 3080 -870
rect 40 -970 3080 -960
rect 40 -1030 3266 -1020
rect 40 -1120 860 -1030
rect 920 -1120 1260 -1030
rect 1320 -1120 1660 -1030
rect 1720 -1120 2790 -1030
rect 2890 -1120 3266 -1030
rect 40 -1130 3266 -1120
<< labels >>
rlabel metal1 2900 850 2900 850 1 net1
port 1 n
rlabel metal1 2940 10 2940 10 1 net3
port 2 n
rlabel metal1 2960 -150 2960 -150 1 net4
port 4 n
rlabel metal1 3010 -1080 3010 -1080 1 net2
port 3 n
rlabel psubdiffcont 1290 1120 1290 1120 1 gnd
port 5 n
<< end >>
