magic
tech sky130A
timestamp 1767864285
<< fence >>
rect -30 0 265 270
<< nwell >>
rect -50 135 285 315
<< nmos >>
rect 15 51 30 93
rect 60 51 75 93
rect 160 51 175 93
rect 205 51 220 93
<< pmos >>
rect 45 160 60 219
rect 90 160 105 219
rect 135 160 150 219
rect 180 160 195 219
<< ndiff >>
rect -12 79 15 93
rect -12 62 -8 79
rect 9 62 15 79
rect -12 51 15 62
rect 30 79 60 93
rect 30 62 36 79
rect 54 62 60 79
rect 30 51 60 62
rect 75 77 102 93
rect 75 60 81 77
rect 98 60 102 77
rect 75 51 102 60
rect 133 79 160 93
rect 133 62 137 79
rect 154 62 160 79
rect 133 51 160 62
rect 175 79 205 93
rect 175 62 181 79
rect 199 62 205 79
rect 175 51 205 62
rect 220 79 247 93
rect 220 62 226 79
rect 243 62 247 79
rect 220 51 247 62
<< pdiff >>
rect 18 211 45 219
rect 18 194 22 211
rect 39 194 45 211
rect 18 160 45 194
rect 60 211 90 219
rect 60 194 66 211
rect 84 194 90 211
rect 60 160 90 194
rect 105 211 135 219
rect 105 194 111 211
rect 129 194 135 211
rect 105 160 135 194
rect 150 211 180 219
rect 150 194 156 211
rect 174 194 180 211
rect 150 160 180 194
rect 195 211 222 219
rect 195 194 201 211
rect 218 194 222 211
rect 195 160 222 194
<< ndiffc >>
rect -8 62 9 79
rect 36 62 54 79
rect 81 60 98 77
rect 137 62 154 79
rect 181 62 199 79
rect 226 62 243 79
<< pdiffc >>
rect 22 194 39 211
rect 66 194 84 211
rect 111 194 129 211
rect 156 194 174 211
rect 201 194 218 211
<< psubdiff >>
rect -30 7 265 24
rect -30 -10 -15 7
rect 2 -10 36 7
rect 54 -10 88 7
rect 105 -10 130 7
rect 147 -10 181 7
rect 199 -10 233 7
rect 250 -10 265 7
rect -30 -24 265 -10
<< nsubdiff >>
rect -30 278 265 295
rect -30 261 15 278
rect 32 261 66 278
rect 84 261 109 278
rect 129 261 156 278
rect 174 261 208 278
rect 225 261 265 278
rect -30 246 265 261
<< psubdiffcont >>
rect -15 -10 2 7
rect 36 -10 54 7
rect 88 -10 105 7
rect 130 -10 147 7
rect 181 -10 199 7
rect 233 -10 250 7
<< nsubdiffcont >>
rect 15 261 32 278
rect 66 261 84 278
rect 109 261 129 278
rect 156 261 174 278
rect 208 261 225 278
<< poly >>
rect 45 219 60 232
rect 90 219 105 232
rect 135 219 150 232
rect 180 219 195 232
rect 45 144 60 160
rect 90 144 105 160
rect 45 136 105 144
rect 45 126 65 136
rect 15 119 65 126
rect 82 119 105 136
rect 15 111 105 119
rect 135 143 150 160
rect 180 143 195 160
rect 135 135 195 143
rect 135 118 158 135
rect 175 125 195 135
rect 175 118 220 125
rect 15 93 30 111
rect 60 93 75 111
rect 135 110 220 118
rect 160 93 175 110
rect 205 93 220 110
rect 15 38 30 51
rect 60 38 75 51
rect 160 38 175 51
rect 205 38 220 51
<< polycont >>
rect 65 119 82 136
rect 158 118 175 135
<< locali >>
rect -30 278 265 295
rect -30 261 15 278
rect 32 261 66 278
rect 84 261 109 278
rect 129 261 156 278
rect 174 261 208 278
rect 225 261 265 278
rect -30 246 265 261
rect 18 211 43 246
rect 18 194 22 211
rect 39 194 43 211
rect 18 160 43 194
rect 62 212 88 219
rect 62 194 65 212
rect 85 194 88 212
rect 62 176 88 194
rect 107 211 133 246
rect 107 194 111 211
rect 129 194 133 211
rect 107 160 133 194
rect 152 212 178 219
rect 152 194 155 212
rect 175 194 178 212
rect 152 161 178 194
rect 197 211 222 246
rect 197 194 201 211
rect 218 194 222 211
rect 197 160 222 194
rect 60 139 90 144
rect 60 119 65 139
rect 82 119 90 139
rect 60 113 90 119
rect 61 111 90 113
rect 150 135 180 143
rect 150 118 158 135
rect 175 118 180 135
rect 150 110 180 118
rect -12 79 13 93
rect -12 62 -8 79
rect 11 62 13 79
rect -12 51 13 62
rect 32 62 36 90
rect 53 79 58 90
rect 54 62 58 79
rect 32 51 58 62
rect 77 85 101 93
rect 77 77 102 85
rect 77 44 81 77
rect 98 44 102 77
rect 133 79 158 93
rect 133 62 137 79
rect 154 62 158 79
rect 133 51 158 62
rect 177 79 203 93
rect 177 62 181 79
rect 199 62 203 79
rect 77 43 102 44
rect 177 24 203 62
rect 222 79 247 93
rect 222 62 224 79
rect 243 62 247 79
rect 222 51 247 62
rect -30 7 265 24
rect -30 -10 -15 7
rect 2 -10 36 7
rect 54 -10 88 7
rect 105 -10 130 7
rect 147 -10 181 7
rect 199 -10 233 7
rect 250 -10 265 7
rect -30 -25 265 -10
<< viali >>
rect 15 261 32 278
rect 66 261 84 278
rect 109 261 129 278
rect 156 261 174 278
rect 208 261 225 278
rect 65 211 85 212
rect 65 194 66 211
rect 66 194 84 211
rect 84 194 85 211
rect 155 211 175 212
rect 155 194 156 211
rect 156 194 174 211
rect 174 194 175 211
rect 65 136 82 139
rect 65 122 82 136
rect 158 118 175 135
rect -6 62 9 79
rect 9 62 11 79
rect 36 79 53 90
rect 36 73 53 79
rect 81 60 98 61
rect 81 44 98 60
rect 137 62 154 79
rect 224 62 226 79
rect 226 62 241 79
rect -15 -10 2 7
rect 36 -10 54 7
rect 88 -10 105 7
rect 130 -10 147 7
rect 181 -10 199 7
rect 233 -10 250 7
<< metal1 >>
rect -30 278 265 295
rect -30 261 15 278
rect 32 261 66 278
rect 84 261 109 278
rect 129 261 156 278
rect 174 261 208 278
rect 225 261 265 278
rect -30 246 265 261
rect 62 219 88 220
rect 152 219 178 220
rect -12 212 178 219
rect -12 194 65 212
rect 85 194 155 212
rect 175 194 178 212
rect -12 185 178 194
rect -12 79 14 185
rect 152 160 178 185
rect 60 139 90 156
rect 60 122 65 139
rect 82 122 90 139
rect 60 112 90 122
rect 150 135 180 143
rect 150 118 158 135
rect 175 118 180 135
rect 150 110 180 118
rect -12 62 -6 79
rect 11 62 14 79
rect 32 90 133 98
rect 32 73 36 90
rect 53 84 133 90
rect 177 84 203 85
rect 53 83 248 84
rect 53 73 58 83
rect 32 66 58 73
rect 119 79 248 83
rect -12 52 14 62
rect 77 61 102 68
rect 77 52 81 61
rect -12 44 81 52
rect 98 44 102 61
rect 119 62 137 79
rect 154 62 224 79
rect 241 62 248 79
rect 119 58 248 62
rect -12 38 102 44
rect -30 7 265 24
rect -30 -10 -15 7
rect 2 -10 36 7
rect 54 -10 88 7
rect 105 -10 130 7
rect 147 -10 181 7
rect 199 -10 233 7
rect 250 -10 265 7
rect -30 -25 265 -10
<< labels >>
rlabel nwell -21 253 254 287 1 vdd
port 1 n
rlabel metal1 -21 -18 254 16 1 gnd
port 2 n
rlabel metal1 155 115 176 133 1 b
port 4 n
rlabel metal1 62 116 88 134 1 a
port 5 n
rlabel metal1 -5 114 8 129 1 out
port 6 n
<< end >>
