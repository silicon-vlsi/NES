magic
tech sky130A
magscale 1 2
timestamp 1764841004
<< pwell >>
rect 0 3850 334 3886
rect 1112 3850 1340 3864
rect 0 3733 1340 3850
rect 0 2699 153 3733
rect 1187 2699 1340 3733
rect 0 2546 1340 2699
rect 1342 3733 2682 3864
rect 1342 2699 1495 3733
rect 2529 2699 2682 3733
rect 1342 2546 2682 2699
rect 2684 3733 4024 3864
rect 2684 2699 2837 3733
rect 3871 2699 4024 3733
rect 2684 2546 4024 2699
rect 4026 3733 5366 3864
rect 4026 2699 4179 3733
rect 5213 2699 5366 3733
rect 4026 2546 5366 2699
rect 5368 3733 6708 3864
rect 5368 2699 5521 3733
rect 6555 2699 6708 3733
rect 5368 2546 6708 2699
rect 6710 3733 8050 3864
rect 6710 2699 6863 3733
rect 7897 2699 8050 3733
rect 6710 2546 8050 2699
rect 8052 3733 9392 3864
rect 8052 2699 8205 3733
rect 9239 2699 9392 3733
rect 8052 2546 9392 2699
rect 0 2391 1340 2544
rect 0 1357 153 2391
rect 1187 1357 1340 2391
rect 0 1204 1340 1357
rect 1342 2391 2682 2544
rect 1342 1357 1495 2391
rect 2529 1357 2682 2391
rect 1342 1204 2682 1357
rect 2684 2391 4024 2544
rect 2684 1357 2837 2391
rect 3871 1357 4024 2391
rect 2684 1204 4024 1357
rect 4026 2391 5366 2544
rect 4026 1357 4179 2391
rect 5213 1357 5366 2391
rect 4026 1204 5366 1357
rect 5368 2391 6708 2544
rect 5368 1357 5521 2391
rect 6555 1357 6708 2391
rect 5368 1204 6708 1357
rect 6710 2391 8050 2544
rect 6710 1357 6863 2391
rect 7897 1357 8050 2391
rect 6710 1204 8050 1357
rect 8052 2391 9392 2544
rect 8052 1357 8205 2391
rect 9239 1357 9392 2391
rect 8052 1204 9392 1357
rect 1686 1049 2682 1177
rect 1342 15 1495 874
rect 2529 15 2682 1049
rect 1342 -138 2682 15
rect 2684 1049 4024 1177
rect 2684 15 2837 1049
rect 3871 15 4024 1049
rect 2684 -138 4024 15
rect 4026 1049 5366 1177
rect 4026 15 4179 1049
rect 5213 15 5366 1049
rect 4026 -138 5366 15
rect 5368 1049 6708 1177
rect 5368 15 5521 1049
rect 6555 15 6708 1049
rect 5368 -138 6708 15
rect 6710 1049 8050 1202
rect 6710 15 6863 1049
rect 7897 15 8050 1049
rect 6710 -138 8050 15
rect 8052 1049 9392 1202
rect 8052 15 8205 1049
rect 9239 15 9392 1049
rect 8052 -138 9392 15
rect 0 -293 1340 -140
rect 0 -1327 153 -293
rect 1187 -1327 1340 -293
rect 0 -1480 1340 -1327
rect 1342 -293 2682 -140
rect 1342 -1327 1495 -293
rect 2529 -1327 2682 -293
rect 1342 -1480 2682 -1327
rect 2684 -293 4024 -140
rect 2684 -1327 2837 -293
rect 3871 -1327 4024 -293
rect 2684 -1480 4024 -1327
rect 4026 -293 5366 -140
rect 4026 -1327 4179 -293
rect 5213 -1327 5366 -293
rect 4026 -1480 5366 -1327
rect 5368 -293 6708 -140
rect 5368 -1327 5521 -293
rect 6555 -1327 6708 -293
rect 5368 -1480 6708 -1327
rect 6710 -293 8050 -140
rect 6710 -1327 6863 -293
rect 7897 -1327 8050 -293
rect 6710 -1480 8050 -1327
rect 8052 -293 9392 -140
rect 8052 -1327 8205 -293
rect 9239 -1327 9392 -293
rect 8052 -1480 9392 -1327
<< nbase >>
rect 153 2699 1187 3733
rect 1495 2699 2529 3733
rect 2837 2699 3871 3733
rect 4179 2699 5213 3733
rect 5521 2699 6555 3733
rect 6863 2699 7897 3733
rect 8205 2699 9239 3733
rect 153 1357 1187 2391
rect 1495 1357 2529 2391
rect 2837 1357 3871 2391
rect 4179 1357 5213 2391
rect 5521 1357 6555 2391
rect 6863 1357 7897 2391
rect 8205 1357 9239 2391
rect 1686 874 2529 1049
rect 1495 15 2529 874
rect 2837 15 3871 1049
rect 4179 15 5213 1049
rect 5521 15 6555 1049
rect 6863 15 7897 1049
rect 8205 15 9239 1049
rect 153 -1327 1187 -293
rect 1495 -1327 2529 -293
rect 2837 -1327 3871 -293
rect 4179 -1327 5213 -293
rect 5521 -1327 6555 -293
rect 6863 -1327 7897 -293
rect 8205 -1327 9239 -293
<< pdiff >>
rect 330 3504 1010 3556
rect 330 3470 384 3504
rect 418 3470 474 3504
rect 508 3470 564 3504
rect 598 3470 654 3504
rect 688 3470 744 3504
rect 778 3470 834 3504
rect 868 3470 924 3504
rect 958 3470 1010 3504
rect 330 3414 1010 3470
rect 330 3380 384 3414
rect 418 3380 474 3414
rect 508 3380 564 3414
rect 598 3380 654 3414
rect 688 3380 744 3414
rect 778 3380 834 3414
rect 868 3380 924 3414
rect 958 3380 1010 3414
rect 330 3324 1010 3380
rect 330 3290 384 3324
rect 418 3290 474 3324
rect 508 3290 564 3324
rect 598 3290 654 3324
rect 688 3290 744 3324
rect 778 3290 834 3324
rect 868 3290 924 3324
rect 958 3290 1010 3324
rect 330 3234 1010 3290
rect 330 3200 384 3234
rect 418 3200 474 3234
rect 508 3200 564 3234
rect 598 3200 654 3234
rect 688 3200 744 3234
rect 778 3200 834 3234
rect 868 3200 924 3234
rect 958 3200 1010 3234
rect 330 3144 1010 3200
rect 330 3110 384 3144
rect 418 3110 474 3144
rect 508 3110 564 3144
rect 598 3110 654 3144
rect 688 3110 744 3144
rect 778 3110 834 3144
rect 868 3110 924 3144
rect 958 3110 1010 3144
rect 330 3054 1010 3110
rect 330 3020 384 3054
rect 418 3020 474 3054
rect 508 3020 564 3054
rect 598 3020 654 3054
rect 688 3020 744 3054
rect 778 3020 834 3054
rect 868 3020 924 3054
rect 958 3020 1010 3054
rect 330 2964 1010 3020
rect 330 2930 384 2964
rect 418 2930 474 2964
rect 508 2930 564 2964
rect 598 2930 654 2964
rect 688 2930 744 2964
rect 778 2930 834 2964
rect 868 2930 924 2964
rect 958 2930 1010 2964
rect 330 2876 1010 2930
rect 1672 3504 2352 3556
rect 1672 3470 1726 3504
rect 1760 3470 1816 3504
rect 1850 3470 1906 3504
rect 1940 3470 1996 3504
rect 2030 3470 2086 3504
rect 2120 3470 2176 3504
rect 2210 3470 2266 3504
rect 2300 3470 2352 3504
rect 1672 3414 2352 3470
rect 1672 3380 1726 3414
rect 1760 3380 1816 3414
rect 1850 3380 1906 3414
rect 1940 3380 1996 3414
rect 2030 3380 2086 3414
rect 2120 3380 2176 3414
rect 2210 3380 2266 3414
rect 2300 3380 2352 3414
rect 1672 3324 2352 3380
rect 1672 3290 1726 3324
rect 1760 3290 1816 3324
rect 1850 3290 1906 3324
rect 1940 3290 1996 3324
rect 2030 3290 2086 3324
rect 2120 3290 2176 3324
rect 2210 3290 2266 3324
rect 2300 3290 2352 3324
rect 1672 3234 2352 3290
rect 1672 3200 1726 3234
rect 1760 3200 1816 3234
rect 1850 3200 1906 3234
rect 1940 3200 1996 3234
rect 2030 3200 2086 3234
rect 2120 3200 2176 3234
rect 2210 3200 2266 3234
rect 2300 3200 2352 3234
rect 1672 3144 2352 3200
rect 1672 3110 1726 3144
rect 1760 3110 1816 3144
rect 1850 3110 1906 3144
rect 1940 3110 1996 3144
rect 2030 3110 2086 3144
rect 2120 3110 2176 3144
rect 2210 3110 2266 3144
rect 2300 3110 2352 3144
rect 1672 3054 2352 3110
rect 1672 3020 1726 3054
rect 1760 3020 1816 3054
rect 1850 3020 1906 3054
rect 1940 3020 1996 3054
rect 2030 3020 2086 3054
rect 2120 3020 2176 3054
rect 2210 3020 2266 3054
rect 2300 3020 2352 3054
rect 1672 2964 2352 3020
rect 1672 2930 1726 2964
rect 1760 2930 1816 2964
rect 1850 2930 1906 2964
rect 1940 2930 1996 2964
rect 2030 2930 2086 2964
rect 2120 2930 2176 2964
rect 2210 2930 2266 2964
rect 2300 2930 2352 2964
rect 1672 2876 2352 2930
rect 3014 3504 3694 3556
rect 3014 3470 3068 3504
rect 3102 3470 3158 3504
rect 3192 3470 3248 3504
rect 3282 3470 3338 3504
rect 3372 3470 3428 3504
rect 3462 3470 3518 3504
rect 3552 3470 3608 3504
rect 3642 3470 3694 3504
rect 3014 3414 3694 3470
rect 3014 3380 3068 3414
rect 3102 3380 3158 3414
rect 3192 3380 3248 3414
rect 3282 3380 3338 3414
rect 3372 3380 3428 3414
rect 3462 3380 3518 3414
rect 3552 3380 3608 3414
rect 3642 3380 3694 3414
rect 3014 3324 3694 3380
rect 3014 3290 3068 3324
rect 3102 3290 3158 3324
rect 3192 3290 3248 3324
rect 3282 3290 3338 3324
rect 3372 3290 3428 3324
rect 3462 3290 3518 3324
rect 3552 3290 3608 3324
rect 3642 3290 3694 3324
rect 3014 3234 3694 3290
rect 3014 3200 3068 3234
rect 3102 3200 3158 3234
rect 3192 3200 3248 3234
rect 3282 3200 3338 3234
rect 3372 3200 3428 3234
rect 3462 3200 3518 3234
rect 3552 3200 3608 3234
rect 3642 3200 3694 3234
rect 3014 3144 3694 3200
rect 3014 3110 3068 3144
rect 3102 3110 3158 3144
rect 3192 3110 3248 3144
rect 3282 3110 3338 3144
rect 3372 3110 3428 3144
rect 3462 3110 3518 3144
rect 3552 3110 3608 3144
rect 3642 3110 3694 3144
rect 3014 3054 3694 3110
rect 3014 3020 3068 3054
rect 3102 3020 3158 3054
rect 3192 3020 3248 3054
rect 3282 3020 3338 3054
rect 3372 3020 3428 3054
rect 3462 3020 3518 3054
rect 3552 3020 3608 3054
rect 3642 3020 3694 3054
rect 3014 2964 3694 3020
rect 3014 2930 3068 2964
rect 3102 2930 3158 2964
rect 3192 2930 3248 2964
rect 3282 2930 3338 2964
rect 3372 2930 3428 2964
rect 3462 2930 3518 2964
rect 3552 2930 3608 2964
rect 3642 2930 3694 2964
rect 3014 2876 3694 2930
rect 4356 3504 5036 3556
rect 4356 3470 4410 3504
rect 4444 3470 4500 3504
rect 4534 3470 4590 3504
rect 4624 3470 4680 3504
rect 4714 3470 4770 3504
rect 4804 3470 4860 3504
rect 4894 3470 4950 3504
rect 4984 3470 5036 3504
rect 4356 3414 5036 3470
rect 4356 3380 4410 3414
rect 4444 3380 4500 3414
rect 4534 3380 4590 3414
rect 4624 3380 4680 3414
rect 4714 3380 4770 3414
rect 4804 3380 4860 3414
rect 4894 3380 4950 3414
rect 4984 3380 5036 3414
rect 4356 3324 5036 3380
rect 4356 3290 4410 3324
rect 4444 3290 4500 3324
rect 4534 3290 4590 3324
rect 4624 3290 4680 3324
rect 4714 3290 4770 3324
rect 4804 3290 4860 3324
rect 4894 3290 4950 3324
rect 4984 3290 5036 3324
rect 4356 3234 5036 3290
rect 4356 3200 4410 3234
rect 4444 3200 4500 3234
rect 4534 3200 4590 3234
rect 4624 3200 4680 3234
rect 4714 3200 4770 3234
rect 4804 3200 4860 3234
rect 4894 3200 4950 3234
rect 4984 3200 5036 3234
rect 4356 3144 5036 3200
rect 4356 3110 4410 3144
rect 4444 3110 4500 3144
rect 4534 3110 4590 3144
rect 4624 3110 4680 3144
rect 4714 3110 4770 3144
rect 4804 3110 4860 3144
rect 4894 3110 4950 3144
rect 4984 3110 5036 3144
rect 4356 3054 5036 3110
rect 4356 3020 4410 3054
rect 4444 3020 4500 3054
rect 4534 3020 4590 3054
rect 4624 3020 4680 3054
rect 4714 3020 4770 3054
rect 4804 3020 4860 3054
rect 4894 3020 4950 3054
rect 4984 3020 5036 3054
rect 4356 2964 5036 3020
rect 4356 2930 4410 2964
rect 4444 2930 4500 2964
rect 4534 2930 4590 2964
rect 4624 2930 4680 2964
rect 4714 2930 4770 2964
rect 4804 2930 4860 2964
rect 4894 2930 4950 2964
rect 4984 2930 5036 2964
rect 4356 2876 5036 2930
rect 5698 3504 6378 3556
rect 5698 3470 5752 3504
rect 5786 3470 5842 3504
rect 5876 3470 5932 3504
rect 5966 3470 6022 3504
rect 6056 3470 6112 3504
rect 6146 3470 6202 3504
rect 6236 3470 6292 3504
rect 6326 3470 6378 3504
rect 5698 3414 6378 3470
rect 5698 3380 5752 3414
rect 5786 3380 5842 3414
rect 5876 3380 5932 3414
rect 5966 3380 6022 3414
rect 6056 3380 6112 3414
rect 6146 3380 6202 3414
rect 6236 3380 6292 3414
rect 6326 3380 6378 3414
rect 5698 3324 6378 3380
rect 5698 3290 5752 3324
rect 5786 3290 5842 3324
rect 5876 3290 5932 3324
rect 5966 3290 6022 3324
rect 6056 3290 6112 3324
rect 6146 3290 6202 3324
rect 6236 3290 6292 3324
rect 6326 3290 6378 3324
rect 5698 3234 6378 3290
rect 5698 3200 5752 3234
rect 5786 3200 5842 3234
rect 5876 3200 5932 3234
rect 5966 3200 6022 3234
rect 6056 3200 6112 3234
rect 6146 3200 6202 3234
rect 6236 3200 6292 3234
rect 6326 3200 6378 3234
rect 5698 3144 6378 3200
rect 5698 3110 5752 3144
rect 5786 3110 5842 3144
rect 5876 3110 5932 3144
rect 5966 3110 6022 3144
rect 6056 3110 6112 3144
rect 6146 3110 6202 3144
rect 6236 3110 6292 3144
rect 6326 3110 6378 3144
rect 5698 3054 6378 3110
rect 5698 3020 5752 3054
rect 5786 3020 5842 3054
rect 5876 3020 5932 3054
rect 5966 3020 6022 3054
rect 6056 3020 6112 3054
rect 6146 3020 6202 3054
rect 6236 3020 6292 3054
rect 6326 3020 6378 3054
rect 5698 2964 6378 3020
rect 5698 2930 5752 2964
rect 5786 2930 5842 2964
rect 5876 2930 5932 2964
rect 5966 2930 6022 2964
rect 6056 2930 6112 2964
rect 6146 2930 6202 2964
rect 6236 2930 6292 2964
rect 6326 2930 6378 2964
rect 5698 2876 6378 2930
rect 7040 3504 7720 3556
rect 7040 3470 7094 3504
rect 7128 3470 7184 3504
rect 7218 3470 7274 3504
rect 7308 3470 7364 3504
rect 7398 3470 7454 3504
rect 7488 3470 7544 3504
rect 7578 3470 7634 3504
rect 7668 3470 7720 3504
rect 7040 3414 7720 3470
rect 7040 3380 7094 3414
rect 7128 3380 7184 3414
rect 7218 3380 7274 3414
rect 7308 3380 7364 3414
rect 7398 3380 7454 3414
rect 7488 3380 7544 3414
rect 7578 3380 7634 3414
rect 7668 3380 7720 3414
rect 7040 3324 7720 3380
rect 7040 3290 7094 3324
rect 7128 3290 7184 3324
rect 7218 3290 7274 3324
rect 7308 3290 7364 3324
rect 7398 3290 7454 3324
rect 7488 3290 7544 3324
rect 7578 3290 7634 3324
rect 7668 3290 7720 3324
rect 7040 3234 7720 3290
rect 7040 3200 7094 3234
rect 7128 3200 7184 3234
rect 7218 3200 7274 3234
rect 7308 3200 7364 3234
rect 7398 3200 7454 3234
rect 7488 3200 7544 3234
rect 7578 3200 7634 3234
rect 7668 3200 7720 3234
rect 7040 3144 7720 3200
rect 7040 3110 7094 3144
rect 7128 3110 7184 3144
rect 7218 3110 7274 3144
rect 7308 3110 7364 3144
rect 7398 3110 7454 3144
rect 7488 3110 7544 3144
rect 7578 3110 7634 3144
rect 7668 3110 7720 3144
rect 7040 3054 7720 3110
rect 7040 3020 7094 3054
rect 7128 3020 7184 3054
rect 7218 3020 7274 3054
rect 7308 3020 7364 3054
rect 7398 3020 7454 3054
rect 7488 3020 7544 3054
rect 7578 3020 7634 3054
rect 7668 3020 7720 3054
rect 7040 2964 7720 3020
rect 7040 2930 7094 2964
rect 7128 2930 7184 2964
rect 7218 2930 7274 2964
rect 7308 2930 7364 2964
rect 7398 2930 7454 2964
rect 7488 2930 7544 2964
rect 7578 2930 7634 2964
rect 7668 2930 7720 2964
rect 7040 2876 7720 2930
rect 8382 3504 9062 3556
rect 8382 3470 8436 3504
rect 8470 3470 8526 3504
rect 8560 3470 8616 3504
rect 8650 3470 8706 3504
rect 8740 3470 8796 3504
rect 8830 3470 8886 3504
rect 8920 3470 8976 3504
rect 9010 3470 9062 3504
rect 8382 3414 9062 3470
rect 8382 3380 8436 3414
rect 8470 3380 8526 3414
rect 8560 3380 8616 3414
rect 8650 3380 8706 3414
rect 8740 3380 8796 3414
rect 8830 3380 8886 3414
rect 8920 3380 8976 3414
rect 9010 3380 9062 3414
rect 8382 3324 9062 3380
rect 8382 3290 8436 3324
rect 8470 3290 8526 3324
rect 8560 3290 8616 3324
rect 8650 3290 8706 3324
rect 8740 3290 8796 3324
rect 8830 3290 8886 3324
rect 8920 3290 8976 3324
rect 9010 3290 9062 3324
rect 8382 3234 9062 3290
rect 8382 3200 8436 3234
rect 8470 3200 8526 3234
rect 8560 3200 8616 3234
rect 8650 3200 8706 3234
rect 8740 3200 8796 3234
rect 8830 3200 8886 3234
rect 8920 3200 8976 3234
rect 9010 3200 9062 3234
rect 8382 3144 9062 3200
rect 8382 3110 8436 3144
rect 8470 3110 8526 3144
rect 8560 3110 8616 3144
rect 8650 3110 8706 3144
rect 8740 3110 8796 3144
rect 8830 3110 8886 3144
rect 8920 3110 8976 3144
rect 9010 3110 9062 3144
rect 8382 3054 9062 3110
rect 8382 3020 8436 3054
rect 8470 3020 8526 3054
rect 8560 3020 8616 3054
rect 8650 3020 8706 3054
rect 8740 3020 8796 3054
rect 8830 3020 8886 3054
rect 8920 3020 8976 3054
rect 9010 3020 9062 3054
rect 8382 2964 9062 3020
rect 8382 2930 8436 2964
rect 8470 2930 8526 2964
rect 8560 2930 8616 2964
rect 8650 2930 8706 2964
rect 8740 2930 8796 2964
rect 8830 2930 8886 2964
rect 8920 2930 8976 2964
rect 9010 2930 9062 2964
rect 8382 2876 9062 2930
rect 330 2162 1010 2214
rect 330 2128 384 2162
rect 418 2128 474 2162
rect 508 2128 564 2162
rect 598 2128 654 2162
rect 688 2128 744 2162
rect 778 2128 834 2162
rect 868 2128 924 2162
rect 958 2128 1010 2162
rect 330 2072 1010 2128
rect 330 2038 384 2072
rect 418 2038 474 2072
rect 508 2038 564 2072
rect 598 2038 654 2072
rect 688 2038 744 2072
rect 778 2038 834 2072
rect 868 2038 924 2072
rect 958 2038 1010 2072
rect 330 1982 1010 2038
rect 330 1948 384 1982
rect 418 1948 474 1982
rect 508 1948 564 1982
rect 598 1948 654 1982
rect 688 1948 744 1982
rect 778 1948 834 1982
rect 868 1948 924 1982
rect 958 1948 1010 1982
rect 330 1892 1010 1948
rect 330 1858 384 1892
rect 418 1858 474 1892
rect 508 1858 564 1892
rect 598 1858 654 1892
rect 688 1858 744 1892
rect 778 1858 834 1892
rect 868 1858 924 1892
rect 958 1858 1010 1892
rect 330 1802 1010 1858
rect 330 1768 384 1802
rect 418 1768 474 1802
rect 508 1768 564 1802
rect 598 1768 654 1802
rect 688 1768 744 1802
rect 778 1768 834 1802
rect 868 1768 924 1802
rect 958 1768 1010 1802
rect 330 1712 1010 1768
rect 330 1678 384 1712
rect 418 1678 474 1712
rect 508 1678 564 1712
rect 598 1678 654 1712
rect 688 1678 744 1712
rect 778 1678 834 1712
rect 868 1678 924 1712
rect 958 1678 1010 1712
rect 330 1622 1010 1678
rect 330 1588 384 1622
rect 418 1588 474 1622
rect 508 1588 564 1622
rect 598 1588 654 1622
rect 688 1588 744 1622
rect 778 1588 834 1622
rect 868 1588 924 1622
rect 958 1588 1010 1622
rect 330 1534 1010 1588
rect 1672 2162 2352 2214
rect 1672 2128 1726 2162
rect 1760 2128 1816 2162
rect 1850 2128 1906 2162
rect 1940 2128 1996 2162
rect 2030 2128 2086 2162
rect 2120 2128 2176 2162
rect 2210 2128 2266 2162
rect 2300 2128 2352 2162
rect 1672 2072 2352 2128
rect 1672 2038 1726 2072
rect 1760 2038 1816 2072
rect 1850 2038 1906 2072
rect 1940 2038 1996 2072
rect 2030 2038 2086 2072
rect 2120 2038 2176 2072
rect 2210 2038 2266 2072
rect 2300 2038 2352 2072
rect 1672 1982 2352 2038
rect 1672 1948 1726 1982
rect 1760 1948 1816 1982
rect 1850 1948 1906 1982
rect 1940 1948 1996 1982
rect 2030 1948 2086 1982
rect 2120 1948 2176 1982
rect 2210 1948 2266 1982
rect 2300 1948 2352 1982
rect 1672 1892 2352 1948
rect 1672 1858 1726 1892
rect 1760 1858 1816 1892
rect 1850 1858 1906 1892
rect 1940 1858 1996 1892
rect 2030 1858 2086 1892
rect 2120 1858 2176 1892
rect 2210 1858 2266 1892
rect 2300 1858 2352 1892
rect 1672 1802 2352 1858
rect 1672 1768 1726 1802
rect 1760 1768 1816 1802
rect 1850 1768 1906 1802
rect 1940 1768 1996 1802
rect 2030 1768 2086 1802
rect 2120 1768 2176 1802
rect 2210 1768 2266 1802
rect 2300 1768 2352 1802
rect 1672 1712 2352 1768
rect 1672 1678 1726 1712
rect 1760 1678 1816 1712
rect 1850 1678 1906 1712
rect 1940 1678 1996 1712
rect 2030 1678 2086 1712
rect 2120 1678 2176 1712
rect 2210 1678 2266 1712
rect 2300 1678 2352 1712
rect 1672 1622 2352 1678
rect 1672 1588 1726 1622
rect 1760 1588 1816 1622
rect 1850 1588 1906 1622
rect 1940 1588 1996 1622
rect 2030 1588 2086 1622
rect 2120 1588 2176 1622
rect 2210 1588 2266 1622
rect 2300 1588 2352 1622
rect 1672 1534 2352 1588
rect 3014 2162 3694 2214
rect 3014 2128 3068 2162
rect 3102 2128 3158 2162
rect 3192 2128 3248 2162
rect 3282 2128 3338 2162
rect 3372 2128 3428 2162
rect 3462 2128 3518 2162
rect 3552 2128 3608 2162
rect 3642 2128 3694 2162
rect 3014 2072 3694 2128
rect 3014 2038 3068 2072
rect 3102 2038 3158 2072
rect 3192 2038 3248 2072
rect 3282 2038 3338 2072
rect 3372 2038 3428 2072
rect 3462 2038 3518 2072
rect 3552 2038 3608 2072
rect 3642 2038 3694 2072
rect 3014 1982 3694 2038
rect 3014 1948 3068 1982
rect 3102 1948 3158 1982
rect 3192 1948 3248 1982
rect 3282 1948 3338 1982
rect 3372 1948 3428 1982
rect 3462 1948 3518 1982
rect 3552 1948 3608 1982
rect 3642 1948 3694 1982
rect 3014 1892 3694 1948
rect 3014 1858 3068 1892
rect 3102 1858 3158 1892
rect 3192 1858 3248 1892
rect 3282 1858 3338 1892
rect 3372 1858 3428 1892
rect 3462 1858 3518 1892
rect 3552 1858 3608 1892
rect 3642 1858 3694 1892
rect 3014 1802 3694 1858
rect 3014 1768 3068 1802
rect 3102 1768 3158 1802
rect 3192 1768 3248 1802
rect 3282 1768 3338 1802
rect 3372 1768 3428 1802
rect 3462 1768 3518 1802
rect 3552 1768 3608 1802
rect 3642 1768 3694 1802
rect 3014 1712 3694 1768
rect 3014 1678 3068 1712
rect 3102 1678 3158 1712
rect 3192 1678 3248 1712
rect 3282 1678 3338 1712
rect 3372 1678 3428 1712
rect 3462 1678 3518 1712
rect 3552 1678 3608 1712
rect 3642 1678 3694 1712
rect 3014 1622 3694 1678
rect 3014 1588 3068 1622
rect 3102 1588 3158 1622
rect 3192 1588 3248 1622
rect 3282 1588 3338 1622
rect 3372 1588 3428 1622
rect 3462 1588 3518 1622
rect 3552 1588 3608 1622
rect 3642 1588 3694 1622
rect 3014 1534 3694 1588
rect 4356 2162 5036 2214
rect 4356 2128 4410 2162
rect 4444 2128 4500 2162
rect 4534 2128 4590 2162
rect 4624 2128 4680 2162
rect 4714 2128 4770 2162
rect 4804 2128 4860 2162
rect 4894 2128 4950 2162
rect 4984 2128 5036 2162
rect 4356 2072 5036 2128
rect 4356 2038 4410 2072
rect 4444 2038 4500 2072
rect 4534 2038 4590 2072
rect 4624 2038 4680 2072
rect 4714 2038 4770 2072
rect 4804 2038 4860 2072
rect 4894 2038 4950 2072
rect 4984 2038 5036 2072
rect 4356 1982 5036 2038
rect 4356 1948 4410 1982
rect 4444 1948 4500 1982
rect 4534 1948 4590 1982
rect 4624 1948 4680 1982
rect 4714 1948 4770 1982
rect 4804 1948 4860 1982
rect 4894 1948 4950 1982
rect 4984 1948 5036 1982
rect 4356 1892 5036 1948
rect 4356 1858 4410 1892
rect 4444 1858 4500 1892
rect 4534 1858 4590 1892
rect 4624 1858 4680 1892
rect 4714 1858 4770 1892
rect 4804 1858 4860 1892
rect 4894 1858 4950 1892
rect 4984 1858 5036 1892
rect 4356 1802 5036 1858
rect 4356 1768 4410 1802
rect 4444 1768 4500 1802
rect 4534 1768 4590 1802
rect 4624 1768 4680 1802
rect 4714 1768 4770 1802
rect 4804 1768 4860 1802
rect 4894 1768 4950 1802
rect 4984 1768 5036 1802
rect 4356 1712 5036 1768
rect 4356 1678 4410 1712
rect 4444 1678 4500 1712
rect 4534 1678 4590 1712
rect 4624 1678 4680 1712
rect 4714 1678 4770 1712
rect 4804 1678 4860 1712
rect 4894 1678 4950 1712
rect 4984 1678 5036 1712
rect 4356 1622 5036 1678
rect 4356 1588 4410 1622
rect 4444 1588 4500 1622
rect 4534 1588 4590 1622
rect 4624 1588 4680 1622
rect 4714 1588 4770 1622
rect 4804 1588 4860 1622
rect 4894 1588 4950 1622
rect 4984 1588 5036 1622
rect 4356 1534 5036 1588
rect 5698 2162 6378 2214
rect 5698 2128 5752 2162
rect 5786 2128 5842 2162
rect 5876 2128 5932 2162
rect 5966 2128 6022 2162
rect 6056 2128 6112 2162
rect 6146 2128 6202 2162
rect 6236 2128 6292 2162
rect 6326 2128 6378 2162
rect 5698 2072 6378 2128
rect 5698 2038 5752 2072
rect 5786 2038 5842 2072
rect 5876 2038 5932 2072
rect 5966 2038 6022 2072
rect 6056 2038 6112 2072
rect 6146 2038 6202 2072
rect 6236 2038 6292 2072
rect 6326 2038 6378 2072
rect 5698 1982 6378 2038
rect 5698 1948 5752 1982
rect 5786 1948 5842 1982
rect 5876 1948 5932 1982
rect 5966 1948 6022 1982
rect 6056 1948 6112 1982
rect 6146 1948 6202 1982
rect 6236 1948 6292 1982
rect 6326 1948 6378 1982
rect 5698 1892 6378 1948
rect 5698 1858 5752 1892
rect 5786 1858 5842 1892
rect 5876 1858 5932 1892
rect 5966 1858 6022 1892
rect 6056 1858 6112 1892
rect 6146 1858 6202 1892
rect 6236 1858 6292 1892
rect 6326 1858 6378 1892
rect 5698 1802 6378 1858
rect 5698 1768 5752 1802
rect 5786 1768 5842 1802
rect 5876 1768 5932 1802
rect 5966 1768 6022 1802
rect 6056 1768 6112 1802
rect 6146 1768 6202 1802
rect 6236 1768 6292 1802
rect 6326 1768 6378 1802
rect 5698 1712 6378 1768
rect 5698 1678 5752 1712
rect 5786 1678 5842 1712
rect 5876 1678 5932 1712
rect 5966 1678 6022 1712
rect 6056 1678 6112 1712
rect 6146 1678 6202 1712
rect 6236 1678 6292 1712
rect 6326 1678 6378 1712
rect 5698 1622 6378 1678
rect 5698 1588 5752 1622
rect 5786 1588 5842 1622
rect 5876 1588 5932 1622
rect 5966 1588 6022 1622
rect 6056 1588 6112 1622
rect 6146 1588 6202 1622
rect 6236 1588 6292 1622
rect 6326 1588 6378 1622
rect 5698 1534 6378 1588
rect 7040 2162 7720 2214
rect 7040 2128 7094 2162
rect 7128 2128 7184 2162
rect 7218 2128 7274 2162
rect 7308 2128 7364 2162
rect 7398 2128 7454 2162
rect 7488 2128 7544 2162
rect 7578 2128 7634 2162
rect 7668 2128 7720 2162
rect 7040 2072 7720 2128
rect 7040 2038 7094 2072
rect 7128 2038 7184 2072
rect 7218 2038 7274 2072
rect 7308 2038 7364 2072
rect 7398 2038 7454 2072
rect 7488 2038 7544 2072
rect 7578 2038 7634 2072
rect 7668 2038 7720 2072
rect 7040 1982 7720 2038
rect 7040 1948 7094 1982
rect 7128 1948 7184 1982
rect 7218 1948 7274 1982
rect 7308 1948 7364 1982
rect 7398 1948 7454 1982
rect 7488 1948 7544 1982
rect 7578 1948 7634 1982
rect 7668 1948 7720 1982
rect 7040 1892 7720 1948
rect 7040 1858 7094 1892
rect 7128 1858 7184 1892
rect 7218 1858 7274 1892
rect 7308 1858 7364 1892
rect 7398 1858 7454 1892
rect 7488 1858 7544 1892
rect 7578 1858 7634 1892
rect 7668 1858 7720 1892
rect 7040 1802 7720 1858
rect 7040 1768 7094 1802
rect 7128 1768 7184 1802
rect 7218 1768 7274 1802
rect 7308 1768 7364 1802
rect 7398 1768 7454 1802
rect 7488 1768 7544 1802
rect 7578 1768 7634 1802
rect 7668 1768 7720 1802
rect 7040 1712 7720 1768
rect 7040 1678 7094 1712
rect 7128 1678 7184 1712
rect 7218 1678 7274 1712
rect 7308 1678 7364 1712
rect 7398 1678 7454 1712
rect 7488 1678 7544 1712
rect 7578 1678 7634 1712
rect 7668 1678 7720 1712
rect 7040 1622 7720 1678
rect 7040 1588 7094 1622
rect 7128 1588 7184 1622
rect 7218 1588 7274 1622
rect 7308 1588 7364 1622
rect 7398 1588 7454 1622
rect 7488 1588 7544 1622
rect 7578 1588 7634 1622
rect 7668 1588 7720 1622
rect 7040 1534 7720 1588
rect 8382 2162 9062 2214
rect 8382 2128 8436 2162
rect 8470 2128 8526 2162
rect 8560 2128 8616 2162
rect 8650 2128 8706 2162
rect 8740 2128 8796 2162
rect 8830 2128 8886 2162
rect 8920 2128 8976 2162
rect 9010 2128 9062 2162
rect 8382 2072 9062 2128
rect 8382 2038 8436 2072
rect 8470 2038 8526 2072
rect 8560 2038 8616 2072
rect 8650 2038 8706 2072
rect 8740 2038 8796 2072
rect 8830 2038 8886 2072
rect 8920 2038 8976 2072
rect 9010 2038 9062 2072
rect 8382 1982 9062 2038
rect 8382 1948 8436 1982
rect 8470 1948 8526 1982
rect 8560 1948 8616 1982
rect 8650 1948 8706 1982
rect 8740 1948 8796 1982
rect 8830 1948 8886 1982
rect 8920 1948 8976 1982
rect 9010 1948 9062 1982
rect 8382 1892 9062 1948
rect 8382 1858 8436 1892
rect 8470 1858 8526 1892
rect 8560 1858 8616 1892
rect 8650 1858 8706 1892
rect 8740 1858 8796 1892
rect 8830 1858 8886 1892
rect 8920 1858 8976 1892
rect 9010 1858 9062 1892
rect 8382 1802 9062 1858
rect 8382 1768 8436 1802
rect 8470 1768 8526 1802
rect 8560 1768 8616 1802
rect 8650 1768 8706 1802
rect 8740 1768 8796 1802
rect 8830 1768 8886 1802
rect 8920 1768 8976 1802
rect 9010 1768 9062 1802
rect 8382 1712 9062 1768
rect 8382 1678 8436 1712
rect 8470 1678 8526 1712
rect 8560 1678 8616 1712
rect 8650 1678 8706 1712
rect 8740 1678 8796 1712
rect 8830 1678 8886 1712
rect 8920 1678 8976 1712
rect 9010 1678 9062 1712
rect 8382 1622 9062 1678
rect 8382 1588 8436 1622
rect 8470 1588 8526 1622
rect 8560 1588 8616 1622
rect 8650 1588 8706 1622
rect 8740 1588 8796 1622
rect 8830 1588 8886 1622
rect 8920 1588 8976 1622
rect 9010 1588 9062 1622
rect 8382 1534 9062 1588
rect 1672 192 2352 872
rect 3014 192 3694 872
rect 4356 192 5036 872
rect 5698 192 6378 872
rect 7040 820 7720 872
rect 7040 786 7094 820
rect 7128 786 7184 820
rect 7218 786 7274 820
rect 7308 786 7364 820
rect 7398 786 7454 820
rect 7488 786 7544 820
rect 7578 786 7634 820
rect 7668 786 7720 820
rect 7040 730 7720 786
rect 7040 696 7094 730
rect 7128 696 7184 730
rect 7218 696 7274 730
rect 7308 696 7364 730
rect 7398 696 7454 730
rect 7488 696 7544 730
rect 7578 696 7634 730
rect 7668 696 7720 730
rect 7040 640 7720 696
rect 7040 606 7094 640
rect 7128 606 7184 640
rect 7218 606 7274 640
rect 7308 606 7364 640
rect 7398 606 7454 640
rect 7488 606 7544 640
rect 7578 606 7634 640
rect 7668 606 7720 640
rect 7040 550 7720 606
rect 7040 516 7094 550
rect 7128 516 7184 550
rect 7218 516 7274 550
rect 7308 516 7364 550
rect 7398 516 7454 550
rect 7488 516 7544 550
rect 7578 516 7634 550
rect 7668 516 7720 550
rect 7040 460 7720 516
rect 7040 426 7094 460
rect 7128 426 7184 460
rect 7218 426 7274 460
rect 7308 426 7364 460
rect 7398 426 7454 460
rect 7488 426 7544 460
rect 7578 426 7634 460
rect 7668 426 7720 460
rect 7040 370 7720 426
rect 7040 336 7094 370
rect 7128 336 7184 370
rect 7218 336 7274 370
rect 7308 336 7364 370
rect 7398 336 7454 370
rect 7488 336 7544 370
rect 7578 336 7634 370
rect 7668 336 7720 370
rect 7040 280 7720 336
rect 7040 246 7094 280
rect 7128 246 7184 280
rect 7218 246 7274 280
rect 7308 246 7364 280
rect 7398 246 7454 280
rect 7488 246 7544 280
rect 7578 246 7634 280
rect 7668 246 7720 280
rect 7040 192 7720 246
rect 8382 820 9062 872
rect 8382 786 8436 820
rect 8470 786 8526 820
rect 8560 786 8616 820
rect 8650 786 8706 820
rect 8740 786 8796 820
rect 8830 786 8886 820
rect 8920 786 8976 820
rect 9010 786 9062 820
rect 8382 730 9062 786
rect 8382 696 8436 730
rect 8470 696 8526 730
rect 8560 696 8616 730
rect 8650 696 8706 730
rect 8740 696 8796 730
rect 8830 696 8886 730
rect 8920 696 8976 730
rect 9010 696 9062 730
rect 8382 640 9062 696
rect 8382 606 8436 640
rect 8470 606 8526 640
rect 8560 606 8616 640
rect 8650 606 8706 640
rect 8740 606 8796 640
rect 8830 606 8886 640
rect 8920 606 8976 640
rect 9010 606 9062 640
rect 8382 550 9062 606
rect 8382 516 8436 550
rect 8470 516 8526 550
rect 8560 516 8616 550
rect 8650 516 8706 550
rect 8740 516 8796 550
rect 8830 516 8886 550
rect 8920 516 8976 550
rect 9010 516 9062 550
rect 8382 460 9062 516
rect 8382 426 8436 460
rect 8470 426 8526 460
rect 8560 426 8616 460
rect 8650 426 8706 460
rect 8740 426 8796 460
rect 8830 426 8886 460
rect 8920 426 8976 460
rect 9010 426 9062 460
rect 8382 370 9062 426
rect 8382 336 8436 370
rect 8470 336 8526 370
rect 8560 336 8616 370
rect 8650 336 8706 370
rect 8740 336 8796 370
rect 8830 336 8886 370
rect 8920 336 8976 370
rect 9010 336 9062 370
rect 8382 280 9062 336
rect 8382 246 8436 280
rect 8470 246 8526 280
rect 8560 246 8616 280
rect 8650 246 8706 280
rect 8740 246 8796 280
rect 8830 246 8886 280
rect 8920 246 8976 280
rect 9010 246 9062 280
rect 8382 192 9062 246
rect 330 -1150 1010 -470
rect 1672 -1150 2352 -470
rect 3014 -1150 3694 -470
rect 4356 -1150 5036 -470
rect 5698 -1150 6378 -470
rect 7040 -522 7720 -470
rect 7040 -556 7094 -522
rect 7128 -556 7184 -522
rect 7218 -556 7274 -522
rect 7308 -556 7364 -522
rect 7398 -556 7454 -522
rect 7488 -556 7544 -522
rect 7578 -556 7634 -522
rect 7668 -556 7720 -522
rect 7040 -612 7720 -556
rect 7040 -646 7094 -612
rect 7128 -646 7184 -612
rect 7218 -646 7274 -612
rect 7308 -646 7364 -612
rect 7398 -646 7454 -612
rect 7488 -646 7544 -612
rect 7578 -646 7634 -612
rect 7668 -646 7720 -612
rect 7040 -702 7720 -646
rect 7040 -736 7094 -702
rect 7128 -736 7184 -702
rect 7218 -736 7274 -702
rect 7308 -736 7364 -702
rect 7398 -736 7454 -702
rect 7488 -736 7544 -702
rect 7578 -736 7634 -702
rect 7668 -736 7720 -702
rect 7040 -792 7720 -736
rect 7040 -826 7094 -792
rect 7128 -826 7184 -792
rect 7218 -826 7274 -792
rect 7308 -826 7364 -792
rect 7398 -826 7454 -792
rect 7488 -826 7544 -792
rect 7578 -826 7634 -792
rect 7668 -826 7720 -792
rect 7040 -882 7720 -826
rect 7040 -916 7094 -882
rect 7128 -916 7184 -882
rect 7218 -916 7274 -882
rect 7308 -916 7364 -882
rect 7398 -916 7454 -882
rect 7488 -916 7544 -882
rect 7578 -916 7634 -882
rect 7668 -916 7720 -882
rect 7040 -972 7720 -916
rect 7040 -1006 7094 -972
rect 7128 -1006 7184 -972
rect 7218 -1006 7274 -972
rect 7308 -1006 7364 -972
rect 7398 -1006 7454 -972
rect 7488 -1006 7544 -972
rect 7578 -1006 7634 -972
rect 7668 -1006 7720 -972
rect 7040 -1062 7720 -1006
rect 7040 -1096 7094 -1062
rect 7128 -1096 7184 -1062
rect 7218 -1096 7274 -1062
rect 7308 -1096 7364 -1062
rect 7398 -1096 7454 -1062
rect 7488 -1096 7544 -1062
rect 7578 -1096 7634 -1062
rect 7668 -1096 7720 -1062
rect 7040 -1150 7720 -1096
rect 8382 -522 9062 -470
rect 8382 -556 8436 -522
rect 8470 -556 8526 -522
rect 8560 -556 8616 -522
rect 8650 -556 8706 -522
rect 8740 -556 8796 -522
rect 8830 -556 8886 -522
rect 8920 -556 8976 -522
rect 9010 -556 9062 -522
rect 8382 -612 9062 -556
rect 8382 -646 8436 -612
rect 8470 -646 8526 -612
rect 8560 -646 8616 -612
rect 8650 -646 8706 -612
rect 8740 -646 8796 -612
rect 8830 -646 8886 -612
rect 8920 -646 8976 -612
rect 9010 -646 9062 -612
rect 8382 -702 9062 -646
rect 8382 -736 8436 -702
rect 8470 -736 8526 -702
rect 8560 -736 8616 -702
rect 8650 -736 8706 -702
rect 8740 -736 8796 -702
rect 8830 -736 8886 -702
rect 8920 -736 8976 -702
rect 9010 -736 9062 -702
rect 8382 -792 9062 -736
rect 8382 -826 8436 -792
rect 8470 -826 8526 -792
rect 8560 -826 8616 -792
rect 8650 -826 8706 -792
rect 8740 -826 8796 -792
rect 8830 -826 8886 -792
rect 8920 -826 8976 -792
rect 9010 -826 9062 -792
rect 8382 -882 9062 -826
rect 8382 -916 8436 -882
rect 8470 -916 8526 -882
rect 8560 -916 8616 -882
rect 8650 -916 8706 -882
rect 8740 -916 8796 -882
rect 8830 -916 8886 -882
rect 8920 -916 8976 -882
rect 9010 -916 9062 -882
rect 8382 -972 9062 -916
rect 8382 -1006 8436 -972
rect 8470 -1006 8526 -972
rect 8560 -1006 8616 -972
rect 8650 -1006 8706 -972
rect 8740 -1006 8796 -972
rect 8830 -1006 8886 -972
rect 8920 -1006 8976 -972
rect 9010 -1006 9062 -972
rect 8382 -1062 9062 -1006
rect 8382 -1096 8436 -1062
rect 8470 -1096 8526 -1062
rect 8560 -1096 8616 -1062
rect 8650 -1096 8706 -1062
rect 8740 -1096 8796 -1062
rect 8830 -1096 8886 -1062
rect 8920 -1096 8976 -1062
rect 9010 -1096 9062 -1062
rect 8382 -1150 9062 -1096
<< pdiffc >>
rect 384 3470 418 3504
rect 474 3470 508 3504
rect 564 3470 598 3504
rect 654 3470 688 3504
rect 744 3470 778 3504
rect 834 3470 868 3504
rect 924 3470 958 3504
rect 384 3380 418 3414
rect 474 3380 508 3414
rect 564 3380 598 3414
rect 654 3380 688 3414
rect 744 3380 778 3414
rect 834 3380 868 3414
rect 924 3380 958 3414
rect 384 3290 418 3324
rect 474 3290 508 3324
rect 564 3290 598 3324
rect 654 3290 688 3324
rect 744 3290 778 3324
rect 834 3290 868 3324
rect 924 3290 958 3324
rect 384 3200 418 3234
rect 474 3200 508 3234
rect 564 3200 598 3234
rect 654 3200 688 3234
rect 744 3200 778 3234
rect 834 3200 868 3234
rect 924 3200 958 3234
rect 384 3110 418 3144
rect 474 3110 508 3144
rect 564 3110 598 3144
rect 654 3110 688 3144
rect 744 3110 778 3144
rect 834 3110 868 3144
rect 924 3110 958 3144
rect 384 3020 418 3054
rect 474 3020 508 3054
rect 564 3020 598 3054
rect 654 3020 688 3054
rect 744 3020 778 3054
rect 834 3020 868 3054
rect 924 3020 958 3054
rect 384 2930 418 2964
rect 474 2930 508 2964
rect 564 2930 598 2964
rect 654 2930 688 2964
rect 744 2930 778 2964
rect 834 2930 868 2964
rect 924 2930 958 2964
rect 1726 3470 1760 3504
rect 1816 3470 1850 3504
rect 1906 3470 1940 3504
rect 1996 3470 2030 3504
rect 2086 3470 2120 3504
rect 2176 3470 2210 3504
rect 2266 3470 2300 3504
rect 1726 3380 1760 3414
rect 1816 3380 1850 3414
rect 1906 3380 1940 3414
rect 1996 3380 2030 3414
rect 2086 3380 2120 3414
rect 2176 3380 2210 3414
rect 2266 3380 2300 3414
rect 1726 3290 1760 3324
rect 1816 3290 1850 3324
rect 1906 3290 1940 3324
rect 1996 3290 2030 3324
rect 2086 3290 2120 3324
rect 2176 3290 2210 3324
rect 2266 3290 2300 3324
rect 1726 3200 1760 3234
rect 1816 3200 1850 3234
rect 1906 3200 1940 3234
rect 1996 3200 2030 3234
rect 2086 3200 2120 3234
rect 2176 3200 2210 3234
rect 2266 3200 2300 3234
rect 1726 3110 1760 3144
rect 1816 3110 1850 3144
rect 1906 3110 1940 3144
rect 1996 3110 2030 3144
rect 2086 3110 2120 3144
rect 2176 3110 2210 3144
rect 2266 3110 2300 3144
rect 1726 3020 1760 3054
rect 1816 3020 1850 3054
rect 1906 3020 1940 3054
rect 1996 3020 2030 3054
rect 2086 3020 2120 3054
rect 2176 3020 2210 3054
rect 2266 3020 2300 3054
rect 1726 2930 1760 2964
rect 1816 2930 1850 2964
rect 1906 2930 1940 2964
rect 1996 2930 2030 2964
rect 2086 2930 2120 2964
rect 2176 2930 2210 2964
rect 2266 2930 2300 2964
rect 3068 3470 3102 3504
rect 3158 3470 3192 3504
rect 3248 3470 3282 3504
rect 3338 3470 3372 3504
rect 3428 3470 3462 3504
rect 3518 3470 3552 3504
rect 3608 3470 3642 3504
rect 3068 3380 3102 3414
rect 3158 3380 3192 3414
rect 3248 3380 3282 3414
rect 3338 3380 3372 3414
rect 3428 3380 3462 3414
rect 3518 3380 3552 3414
rect 3608 3380 3642 3414
rect 3068 3290 3102 3324
rect 3158 3290 3192 3324
rect 3248 3290 3282 3324
rect 3338 3290 3372 3324
rect 3428 3290 3462 3324
rect 3518 3290 3552 3324
rect 3608 3290 3642 3324
rect 3068 3200 3102 3234
rect 3158 3200 3192 3234
rect 3248 3200 3282 3234
rect 3338 3200 3372 3234
rect 3428 3200 3462 3234
rect 3518 3200 3552 3234
rect 3608 3200 3642 3234
rect 3068 3110 3102 3144
rect 3158 3110 3192 3144
rect 3248 3110 3282 3144
rect 3338 3110 3372 3144
rect 3428 3110 3462 3144
rect 3518 3110 3552 3144
rect 3608 3110 3642 3144
rect 3068 3020 3102 3054
rect 3158 3020 3192 3054
rect 3248 3020 3282 3054
rect 3338 3020 3372 3054
rect 3428 3020 3462 3054
rect 3518 3020 3552 3054
rect 3608 3020 3642 3054
rect 3068 2930 3102 2964
rect 3158 2930 3192 2964
rect 3248 2930 3282 2964
rect 3338 2930 3372 2964
rect 3428 2930 3462 2964
rect 3518 2930 3552 2964
rect 3608 2930 3642 2964
rect 4410 3470 4444 3504
rect 4500 3470 4534 3504
rect 4590 3470 4624 3504
rect 4680 3470 4714 3504
rect 4770 3470 4804 3504
rect 4860 3470 4894 3504
rect 4950 3470 4984 3504
rect 4410 3380 4444 3414
rect 4500 3380 4534 3414
rect 4590 3380 4624 3414
rect 4680 3380 4714 3414
rect 4770 3380 4804 3414
rect 4860 3380 4894 3414
rect 4950 3380 4984 3414
rect 4410 3290 4444 3324
rect 4500 3290 4534 3324
rect 4590 3290 4624 3324
rect 4680 3290 4714 3324
rect 4770 3290 4804 3324
rect 4860 3290 4894 3324
rect 4950 3290 4984 3324
rect 4410 3200 4444 3234
rect 4500 3200 4534 3234
rect 4590 3200 4624 3234
rect 4680 3200 4714 3234
rect 4770 3200 4804 3234
rect 4860 3200 4894 3234
rect 4950 3200 4984 3234
rect 4410 3110 4444 3144
rect 4500 3110 4534 3144
rect 4590 3110 4624 3144
rect 4680 3110 4714 3144
rect 4770 3110 4804 3144
rect 4860 3110 4894 3144
rect 4950 3110 4984 3144
rect 4410 3020 4444 3054
rect 4500 3020 4534 3054
rect 4590 3020 4624 3054
rect 4680 3020 4714 3054
rect 4770 3020 4804 3054
rect 4860 3020 4894 3054
rect 4950 3020 4984 3054
rect 4410 2930 4444 2964
rect 4500 2930 4534 2964
rect 4590 2930 4624 2964
rect 4680 2930 4714 2964
rect 4770 2930 4804 2964
rect 4860 2930 4894 2964
rect 4950 2930 4984 2964
rect 5752 3470 5786 3504
rect 5842 3470 5876 3504
rect 5932 3470 5966 3504
rect 6022 3470 6056 3504
rect 6112 3470 6146 3504
rect 6202 3470 6236 3504
rect 6292 3470 6326 3504
rect 5752 3380 5786 3414
rect 5842 3380 5876 3414
rect 5932 3380 5966 3414
rect 6022 3380 6056 3414
rect 6112 3380 6146 3414
rect 6202 3380 6236 3414
rect 6292 3380 6326 3414
rect 5752 3290 5786 3324
rect 5842 3290 5876 3324
rect 5932 3290 5966 3324
rect 6022 3290 6056 3324
rect 6112 3290 6146 3324
rect 6202 3290 6236 3324
rect 6292 3290 6326 3324
rect 5752 3200 5786 3234
rect 5842 3200 5876 3234
rect 5932 3200 5966 3234
rect 6022 3200 6056 3234
rect 6112 3200 6146 3234
rect 6202 3200 6236 3234
rect 6292 3200 6326 3234
rect 5752 3110 5786 3144
rect 5842 3110 5876 3144
rect 5932 3110 5966 3144
rect 6022 3110 6056 3144
rect 6112 3110 6146 3144
rect 6202 3110 6236 3144
rect 6292 3110 6326 3144
rect 5752 3020 5786 3054
rect 5842 3020 5876 3054
rect 5932 3020 5966 3054
rect 6022 3020 6056 3054
rect 6112 3020 6146 3054
rect 6202 3020 6236 3054
rect 6292 3020 6326 3054
rect 5752 2930 5786 2964
rect 5842 2930 5876 2964
rect 5932 2930 5966 2964
rect 6022 2930 6056 2964
rect 6112 2930 6146 2964
rect 6202 2930 6236 2964
rect 6292 2930 6326 2964
rect 7094 3470 7128 3504
rect 7184 3470 7218 3504
rect 7274 3470 7308 3504
rect 7364 3470 7398 3504
rect 7454 3470 7488 3504
rect 7544 3470 7578 3504
rect 7634 3470 7668 3504
rect 7094 3380 7128 3414
rect 7184 3380 7218 3414
rect 7274 3380 7308 3414
rect 7364 3380 7398 3414
rect 7454 3380 7488 3414
rect 7544 3380 7578 3414
rect 7634 3380 7668 3414
rect 7094 3290 7128 3324
rect 7184 3290 7218 3324
rect 7274 3290 7308 3324
rect 7364 3290 7398 3324
rect 7454 3290 7488 3324
rect 7544 3290 7578 3324
rect 7634 3290 7668 3324
rect 7094 3200 7128 3234
rect 7184 3200 7218 3234
rect 7274 3200 7308 3234
rect 7364 3200 7398 3234
rect 7454 3200 7488 3234
rect 7544 3200 7578 3234
rect 7634 3200 7668 3234
rect 7094 3110 7128 3144
rect 7184 3110 7218 3144
rect 7274 3110 7308 3144
rect 7364 3110 7398 3144
rect 7454 3110 7488 3144
rect 7544 3110 7578 3144
rect 7634 3110 7668 3144
rect 7094 3020 7128 3054
rect 7184 3020 7218 3054
rect 7274 3020 7308 3054
rect 7364 3020 7398 3054
rect 7454 3020 7488 3054
rect 7544 3020 7578 3054
rect 7634 3020 7668 3054
rect 7094 2930 7128 2964
rect 7184 2930 7218 2964
rect 7274 2930 7308 2964
rect 7364 2930 7398 2964
rect 7454 2930 7488 2964
rect 7544 2930 7578 2964
rect 7634 2930 7668 2964
rect 8436 3470 8470 3504
rect 8526 3470 8560 3504
rect 8616 3470 8650 3504
rect 8706 3470 8740 3504
rect 8796 3470 8830 3504
rect 8886 3470 8920 3504
rect 8976 3470 9010 3504
rect 8436 3380 8470 3414
rect 8526 3380 8560 3414
rect 8616 3380 8650 3414
rect 8706 3380 8740 3414
rect 8796 3380 8830 3414
rect 8886 3380 8920 3414
rect 8976 3380 9010 3414
rect 8436 3290 8470 3324
rect 8526 3290 8560 3324
rect 8616 3290 8650 3324
rect 8706 3290 8740 3324
rect 8796 3290 8830 3324
rect 8886 3290 8920 3324
rect 8976 3290 9010 3324
rect 8436 3200 8470 3234
rect 8526 3200 8560 3234
rect 8616 3200 8650 3234
rect 8706 3200 8740 3234
rect 8796 3200 8830 3234
rect 8886 3200 8920 3234
rect 8976 3200 9010 3234
rect 8436 3110 8470 3144
rect 8526 3110 8560 3144
rect 8616 3110 8650 3144
rect 8706 3110 8740 3144
rect 8796 3110 8830 3144
rect 8886 3110 8920 3144
rect 8976 3110 9010 3144
rect 8436 3020 8470 3054
rect 8526 3020 8560 3054
rect 8616 3020 8650 3054
rect 8706 3020 8740 3054
rect 8796 3020 8830 3054
rect 8886 3020 8920 3054
rect 8976 3020 9010 3054
rect 8436 2930 8470 2964
rect 8526 2930 8560 2964
rect 8616 2930 8650 2964
rect 8706 2930 8740 2964
rect 8796 2930 8830 2964
rect 8886 2930 8920 2964
rect 8976 2930 9010 2964
rect 384 2128 418 2162
rect 474 2128 508 2162
rect 564 2128 598 2162
rect 654 2128 688 2162
rect 744 2128 778 2162
rect 834 2128 868 2162
rect 924 2128 958 2162
rect 384 2038 418 2072
rect 474 2038 508 2072
rect 564 2038 598 2072
rect 654 2038 688 2072
rect 744 2038 778 2072
rect 834 2038 868 2072
rect 924 2038 958 2072
rect 384 1948 418 1982
rect 474 1948 508 1982
rect 564 1948 598 1982
rect 654 1948 688 1982
rect 744 1948 778 1982
rect 834 1948 868 1982
rect 924 1948 958 1982
rect 384 1858 418 1892
rect 474 1858 508 1892
rect 564 1858 598 1892
rect 654 1858 688 1892
rect 744 1858 778 1892
rect 834 1858 868 1892
rect 924 1858 958 1892
rect 384 1768 418 1802
rect 474 1768 508 1802
rect 564 1768 598 1802
rect 654 1768 688 1802
rect 744 1768 778 1802
rect 834 1768 868 1802
rect 924 1768 958 1802
rect 384 1678 418 1712
rect 474 1678 508 1712
rect 564 1678 598 1712
rect 654 1678 688 1712
rect 744 1678 778 1712
rect 834 1678 868 1712
rect 924 1678 958 1712
rect 384 1588 418 1622
rect 474 1588 508 1622
rect 564 1588 598 1622
rect 654 1588 688 1622
rect 744 1588 778 1622
rect 834 1588 868 1622
rect 924 1588 958 1622
rect 1726 2128 1760 2162
rect 1816 2128 1850 2162
rect 1906 2128 1940 2162
rect 1996 2128 2030 2162
rect 2086 2128 2120 2162
rect 2176 2128 2210 2162
rect 2266 2128 2300 2162
rect 1726 2038 1760 2072
rect 1816 2038 1850 2072
rect 1906 2038 1940 2072
rect 1996 2038 2030 2072
rect 2086 2038 2120 2072
rect 2176 2038 2210 2072
rect 2266 2038 2300 2072
rect 1726 1948 1760 1982
rect 1816 1948 1850 1982
rect 1906 1948 1940 1982
rect 1996 1948 2030 1982
rect 2086 1948 2120 1982
rect 2176 1948 2210 1982
rect 2266 1948 2300 1982
rect 1726 1858 1760 1892
rect 1816 1858 1850 1892
rect 1906 1858 1940 1892
rect 1996 1858 2030 1892
rect 2086 1858 2120 1892
rect 2176 1858 2210 1892
rect 2266 1858 2300 1892
rect 1726 1768 1760 1802
rect 1816 1768 1850 1802
rect 1906 1768 1940 1802
rect 1996 1768 2030 1802
rect 2086 1768 2120 1802
rect 2176 1768 2210 1802
rect 2266 1768 2300 1802
rect 1726 1678 1760 1712
rect 1816 1678 1850 1712
rect 1906 1678 1940 1712
rect 1996 1678 2030 1712
rect 2086 1678 2120 1712
rect 2176 1678 2210 1712
rect 2266 1678 2300 1712
rect 1726 1588 1760 1622
rect 1816 1588 1850 1622
rect 1906 1588 1940 1622
rect 1996 1588 2030 1622
rect 2086 1588 2120 1622
rect 2176 1588 2210 1622
rect 2266 1588 2300 1622
rect 3068 2128 3102 2162
rect 3158 2128 3192 2162
rect 3248 2128 3282 2162
rect 3338 2128 3372 2162
rect 3428 2128 3462 2162
rect 3518 2128 3552 2162
rect 3608 2128 3642 2162
rect 3068 2038 3102 2072
rect 3158 2038 3192 2072
rect 3248 2038 3282 2072
rect 3338 2038 3372 2072
rect 3428 2038 3462 2072
rect 3518 2038 3552 2072
rect 3608 2038 3642 2072
rect 3068 1948 3102 1982
rect 3158 1948 3192 1982
rect 3248 1948 3282 1982
rect 3338 1948 3372 1982
rect 3428 1948 3462 1982
rect 3518 1948 3552 1982
rect 3608 1948 3642 1982
rect 3068 1858 3102 1892
rect 3158 1858 3192 1892
rect 3248 1858 3282 1892
rect 3338 1858 3372 1892
rect 3428 1858 3462 1892
rect 3518 1858 3552 1892
rect 3608 1858 3642 1892
rect 3068 1768 3102 1802
rect 3158 1768 3192 1802
rect 3248 1768 3282 1802
rect 3338 1768 3372 1802
rect 3428 1768 3462 1802
rect 3518 1768 3552 1802
rect 3608 1768 3642 1802
rect 3068 1678 3102 1712
rect 3158 1678 3192 1712
rect 3248 1678 3282 1712
rect 3338 1678 3372 1712
rect 3428 1678 3462 1712
rect 3518 1678 3552 1712
rect 3608 1678 3642 1712
rect 3068 1588 3102 1622
rect 3158 1588 3192 1622
rect 3248 1588 3282 1622
rect 3338 1588 3372 1622
rect 3428 1588 3462 1622
rect 3518 1588 3552 1622
rect 3608 1588 3642 1622
rect 4410 2128 4444 2162
rect 4500 2128 4534 2162
rect 4590 2128 4624 2162
rect 4680 2128 4714 2162
rect 4770 2128 4804 2162
rect 4860 2128 4894 2162
rect 4950 2128 4984 2162
rect 4410 2038 4444 2072
rect 4500 2038 4534 2072
rect 4590 2038 4624 2072
rect 4680 2038 4714 2072
rect 4770 2038 4804 2072
rect 4860 2038 4894 2072
rect 4950 2038 4984 2072
rect 4410 1948 4444 1982
rect 4500 1948 4534 1982
rect 4590 1948 4624 1982
rect 4680 1948 4714 1982
rect 4770 1948 4804 1982
rect 4860 1948 4894 1982
rect 4950 1948 4984 1982
rect 4410 1858 4444 1892
rect 4500 1858 4534 1892
rect 4590 1858 4624 1892
rect 4680 1858 4714 1892
rect 4770 1858 4804 1892
rect 4860 1858 4894 1892
rect 4950 1858 4984 1892
rect 4410 1768 4444 1802
rect 4500 1768 4534 1802
rect 4590 1768 4624 1802
rect 4680 1768 4714 1802
rect 4770 1768 4804 1802
rect 4860 1768 4894 1802
rect 4950 1768 4984 1802
rect 4410 1678 4444 1712
rect 4500 1678 4534 1712
rect 4590 1678 4624 1712
rect 4680 1678 4714 1712
rect 4770 1678 4804 1712
rect 4860 1678 4894 1712
rect 4950 1678 4984 1712
rect 4410 1588 4444 1622
rect 4500 1588 4534 1622
rect 4590 1588 4624 1622
rect 4680 1588 4714 1622
rect 4770 1588 4804 1622
rect 4860 1588 4894 1622
rect 4950 1588 4984 1622
rect 5752 2128 5786 2162
rect 5842 2128 5876 2162
rect 5932 2128 5966 2162
rect 6022 2128 6056 2162
rect 6112 2128 6146 2162
rect 6202 2128 6236 2162
rect 6292 2128 6326 2162
rect 5752 2038 5786 2072
rect 5842 2038 5876 2072
rect 5932 2038 5966 2072
rect 6022 2038 6056 2072
rect 6112 2038 6146 2072
rect 6202 2038 6236 2072
rect 6292 2038 6326 2072
rect 5752 1948 5786 1982
rect 5842 1948 5876 1982
rect 5932 1948 5966 1982
rect 6022 1948 6056 1982
rect 6112 1948 6146 1982
rect 6202 1948 6236 1982
rect 6292 1948 6326 1982
rect 5752 1858 5786 1892
rect 5842 1858 5876 1892
rect 5932 1858 5966 1892
rect 6022 1858 6056 1892
rect 6112 1858 6146 1892
rect 6202 1858 6236 1892
rect 6292 1858 6326 1892
rect 5752 1768 5786 1802
rect 5842 1768 5876 1802
rect 5932 1768 5966 1802
rect 6022 1768 6056 1802
rect 6112 1768 6146 1802
rect 6202 1768 6236 1802
rect 6292 1768 6326 1802
rect 5752 1678 5786 1712
rect 5842 1678 5876 1712
rect 5932 1678 5966 1712
rect 6022 1678 6056 1712
rect 6112 1678 6146 1712
rect 6202 1678 6236 1712
rect 6292 1678 6326 1712
rect 5752 1588 5786 1622
rect 5842 1588 5876 1622
rect 5932 1588 5966 1622
rect 6022 1588 6056 1622
rect 6112 1588 6146 1622
rect 6202 1588 6236 1622
rect 6292 1588 6326 1622
rect 7094 2128 7128 2162
rect 7184 2128 7218 2162
rect 7274 2128 7308 2162
rect 7364 2128 7398 2162
rect 7454 2128 7488 2162
rect 7544 2128 7578 2162
rect 7634 2128 7668 2162
rect 7094 2038 7128 2072
rect 7184 2038 7218 2072
rect 7274 2038 7308 2072
rect 7364 2038 7398 2072
rect 7454 2038 7488 2072
rect 7544 2038 7578 2072
rect 7634 2038 7668 2072
rect 7094 1948 7128 1982
rect 7184 1948 7218 1982
rect 7274 1948 7308 1982
rect 7364 1948 7398 1982
rect 7454 1948 7488 1982
rect 7544 1948 7578 1982
rect 7634 1948 7668 1982
rect 7094 1858 7128 1892
rect 7184 1858 7218 1892
rect 7274 1858 7308 1892
rect 7364 1858 7398 1892
rect 7454 1858 7488 1892
rect 7544 1858 7578 1892
rect 7634 1858 7668 1892
rect 7094 1768 7128 1802
rect 7184 1768 7218 1802
rect 7274 1768 7308 1802
rect 7364 1768 7398 1802
rect 7454 1768 7488 1802
rect 7544 1768 7578 1802
rect 7634 1768 7668 1802
rect 7094 1678 7128 1712
rect 7184 1678 7218 1712
rect 7274 1678 7308 1712
rect 7364 1678 7398 1712
rect 7454 1678 7488 1712
rect 7544 1678 7578 1712
rect 7634 1678 7668 1712
rect 7094 1588 7128 1622
rect 7184 1588 7218 1622
rect 7274 1588 7308 1622
rect 7364 1588 7398 1622
rect 7454 1588 7488 1622
rect 7544 1588 7578 1622
rect 7634 1588 7668 1622
rect 8436 2128 8470 2162
rect 8526 2128 8560 2162
rect 8616 2128 8650 2162
rect 8706 2128 8740 2162
rect 8796 2128 8830 2162
rect 8886 2128 8920 2162
rect 8976 2128 9010 2162
rect 8436 2038 8470 2072
rect 8526 2038 8560 2072
rect 8616 2038 8650 2072
rect 8706 2038 8740 2072
rect 8796 2038 8830 2072
rect 8886 2038 8920 2072
rect 8976 2038 9010 2072
rect 8436 1948 8470 1982
rect 8526 1948 8560 1982
rect 8616 1948 8650 1982
rect 8706 1948 8740 1982
rect 8796 1948 8830 1982
rect 8886 1948 8920 1982
rect 8976 1948 9010 1982
rect 8436 1858 8470 1892
rect 8526 1858 8560 1892
rect 8616 1858 8650 1892
rect 8706 1858 8740 1892
rect 8796 1858 8830 1892
rect 8886 1858 8920 1892
rect 8976 1858 9010 1892
rect 8436 1768 8470 1802
rect 8526 1768 8560 1802
rect 8616 1768 8650 1802
rect 8706 1768 8740 1802
rect 8796 1768 8830 1802
rect 8886 1768 8920 1802
rect 8976 1768 9010 1802
rect 8436 1678 8470 1712
rect 8526 1678 8560 1712
rect 8616 1678 8650 1712
rect 8706 1678 8740 1712
rect 8796 1678 8830 1712
rect 8886 1678 8920 1712
rect 8976 1678 9010 1712
rect 8436 1588 8470 1622
rect 8526 1588 8560 1622
rect 8616 1588 8650 1622
rect 8706 1588 8740 1622
rect 8796 1588 8830 1622
rect 8886 1588 8920 1622
rect 8976 1588 9010 1622
rect 7094 786 7128 820
rect 7184 786 7218 820
rect 7274 786 7308 820
rect 7364 786 7398 820
rect 7454 786 7488 820
rect 7544 786 7578 820
rect 7634 786 7668 820
rect 7094 696 7128 730
rect 7184 696 7218 730
rect 7274 696 7308 730
rect 7364 696 7398 730
rect 7454 696 7488 730
rect 7544 696 7578 730
rect 7634 696 7668 730
rect 7094 606 7128 640
rect 7184 606 7218 640
rect 7274 606 7308 640
rect 7364 606 7398 640
rect 7454 606 7488 640
rect 7544 606 7578 640
rect 7634 606 7668 640
rect 7094 516 7128 550
rect 7184 516 7218 550
rect 7274 516 7308 550
rect 7364 516 7398 550
rect 7454 516 7488 550
rect 7544 516 7578 550
rect 7634 516 7668 550
rect 7094 426 7128 460
rect 7184 426 7218 460
rect 7274 426 7308 460
rect 7364 426 7398 460
rect 7454 426 7488 460
rect 7544 426 7578 460
rect 7634 426 7668 460
rect 7094 336 7128 370
rect 7184 336 7218 370
rect 7274 336 7308 370
rect 7364 336 7398 370
rect 7454 336 7488 370
rect 7544 336 7578 370
rect 7634 336 7668 370
rect 7094 246 7128 280
rect 7184 246 7218 280
rect 7274 246 7308 280
rect 7364 246 7398 280
rect 7454 246 7488 280
rect 7544 246 7578 280
rect 7634 246 7668 280
rect 8436 786 8470 820
rect 8526 786 8560 820
rect 8616 786 8650 820
rect 8706 786 8740 820
rect 8796 786 8830 820
rect 8886 786 8920 820
rect 8976 786 9010 820
rect 8436 696 8470 730
rect 8526 696 8560 730
rect 8616 696 8650 730
rect 8706 696 8740 730
rect 8796 696 8830 730
rect 8886 696 8920 730
rect 8976 696 9010 730
rect 8436 606 8470 640
rect 8526 606 8560 640
rect 8616 606 8650 640
rect 8706 606 8740 640
rect 8796 606 8830 640
rect 8886 606 8920 640
rect 8976 606 9010 640
rect 8436 516 8470 550
rect 8526 516 8560 550
rect 8616 516 8650 550
rect 8706 516 8740 550
rect 8796 516 8830 550
rect 8886 516 8920 550
rect 8976 516 9010 550
rect 8436 426 8470 460
rect 8526 426 8560 460
rect 8616 426 8650 460
rect 8706 426 8740 460
rect 8796 426 8830 460
rect 8886 426 8920 460
rect 8976 426 9010 460
rect 8436 336 8470 370
rect 8526 336 8560 370
rect 8616 336 8650 370
rect 8706 336 8740 370
rect 8796 336 8830 370
rect 8886 336 8920 370
rect 8976 336 9010 370
rect 8436 246 8470 280
rect 8526 246 8560 280
rect 8616 246 8650 280
rect 8706 246 8740 280
rect 8796 246 8830 280
rect 8886 246 8920 280
rect 8976 246 9010 280
rect 7094 -556 7128 -522
rect 7184 -556 7218 -522
rect 7274 -556 7308 -522
rect 7364 -556 7398 -522
rect 7454 -556 7488 -522
rect 7544 -556 7578 -522
rect 7634 -556 7668 -522
rect 7094 -646 7128 -612
rect 7184 -646 7218 -612
rect 7274 -646 7308 -612
rect 7364 -646 7398 -612
rect 7454 -646 7488 -612
rect 7544 -646 7578 -612
rect 7634 -646 7668 -612
rect 7094 -736 7128 -702
rect 7184 -736 7218 -702
rect 7274 -736 7308 -702
rect 7364 -736 7398 -702
rect 7454 -736 7488 -702
rect 7544 -736 7578 -702
rect 7634 -736 7668 -702
rect 7094 -826 7128 -792
rect 7184 -826 7218 -792
rect 7274 -826 7308 -792
rect 7364 -826 7398 -792
rect 7454 -826 7488 -792
rect 7544 -826 7578 -792
rect 7634 -826 7668 -792
rect 7094 -916 7128 -882
rect 7184 -916 7218 -882
rect 7274 -916 7308 -882
rect 7364 -916 7398 -882
rect 7454 -916 7488 -882
rect 7544 -916 7578 -882
rect 7634 -916 7668 -882
rect 7094 -1006 7128 -972
rect 7184 -1006 7218 -972
rect 7274 -1006 7308 -972
rect 7364 -1006 7398 -972
rect 7454 -1006 7488 -972
rect 7544 -1006 7578 -972
rect 7634 -1006 7668 -972
rect 7094 -1096 7128 -1062
rect 7184 -1096 7218 -1062
rect 7274 -1096 7308 -1062
rect 7364 -1096 7398 -1062
rect 7454 -1096 7488 -1062
rect 7544 -1096 7578 -1062
rect 7634 -1096 7668 -1062
rect 8436 -556 8470 -522
rect 8526 -556 8560 -522
rect 8616 -556 8650 -522
rect 8706 -556 8740 -522
rect 8796 -556 8830 -522
rect 8886 -556 8920 -522
rect 8976 -556 9010 -522
rect 8436 -646 8470 -612
rect 8526 -646 8560 -612
rect 8616 -646 8650 -612
rect 8706 -646 8740 -612
rect 8796 -646 8830 -612
rect 8886 -646 8920 -612
rect 8976 -646 9010 -612
rect 8436 -736 8470 -702
rect 8526 -736 8560 -702
rect 8616 -736 8650 -702
rect 8706 -736 8740 -702
rect 8796 -736 8830 -702
rect 8886 -736 8920 -702
rect 8976 -736 9010 -702
rect 8436 -826 8470 -792
rect 8526 -826 8560 -792
rect 8616 -826 8650 -792
rect 8706 -826 8740 -792
rect 8796 -826 8830 -792
rect 8886 -826 8920 -792
rect 8976 -826 9010 -792
rect 8436 -916 8470 -882
rect 8526 -916 8560 -882
rect 8616 -916 8650 -882
rect 8706 -916 8740 -882
rect 8796 -916 8830 -882
rect 8886 -916 8920 -882
rect 8976 -916 9010 -882
rect 8436 -1006 8470 -972
rect 8526 -1006 8560 -972
rect 8616 -1006 8650 -972
rect 8706 -1006 8740 -972
rect 8796 -1006 8830 -972
rect 8886 -1006 8920 -972
rect 8976 -1006 9010 -972
rect 8436 -1096 8470 -1062
rect 8526 -1096 8560 -1062
rect 8616 -1096 8650 -1062
rect 8706 -1096 8740 -1062
rect 8796 -1096 8830 -1062
rect 8886 -1096 8920 -1062
rect 8976 -1096 9010 -1062
<< psubdiff >>
rect 26 3850 334 3860
rect 1112 3850 1314 3860
rect 26 3825 1314 3850
rect 26 3802 156 3825
rect 26 3768 60 3802
rect 94 3791 156 3802
rect 190 3791 246 3825
rect 280 3791 336 3825
rect 370 3791 426 3825
rect 460 3791 516 3825
rect 550 3791 606 3825
rect 640 3791 696 3825
rect 730 3791 786 3825
rect 820 3791 876 3825
rect 910 3791 966 3825
rect 1000 3791 1056 3825
rect 1090 3791 1146 3825
rect 1180 3802 1314 3825
rect 1180 3791 1247 3802
rect 94 3768 1247 3791
rect 1281 3768 1314 3802
rect 26 3759 1314 3768
rect 26 3712 127 3759
rect 26 3678 60 3712
rect 94 3678 127 3712
rect 1213 3712 1314 3759
rect 26 3622 127 3678
rect 26 3588 60 3622
rect 94 3588 127 3622
rect 26 3532 127 3588
rect 26 3498 60 3532
rect 94 3498 127 3532
rect 26 3442 127 3498
rect 26 3408 60 3442
rect 94 3408 127 3442
rect 26 3352 127 3408
rect 26 3318 60 3352
rect 94 3318 127 3352
rect 26 3262 127 3318
rect 26 3228 60 3262
rect 94 3228 127 3262
rect 26 3172 127 3228
rect 26 3138 60 3172
rect 94 3138 127 3172
rect 26 3082 127 3138
rect 26 3048 60 3082
rect 94 3048 127 3082
rect 26 2992 127 3048
rect 26 2958 60 2992
rect 94 2958 127 2992
rect 26 2902 127 2958
rect 26 2868 60 2902
rect 94 2868 127 2902
rect 26 2812 127 2868
rect 26 2778 60 2812
rect 94 2778 127 2812
rect 26 2722 127 2778
rect 1213 3678 1247 3712
rect 1281 3678 1314 3712
rect 1213 3622 1314 3678
rect 1213 3588 1247 3622
rect 1281 3588 1314 3622
rect 1213 3532 1314 3588
rect 1213 3498 1247 3532
rect 1281 3498 1314 3532
rect 1213 3442 1314 3498
rect 1213 3408 1247 3442
rect 1281 3408 1314 3442
rect 1213 3352 1314 3408
rect 1213 3318 1247 3352
rect 1281 3318 1314 3352
rect 1213 3262 1314 3318
rect 1213 3228 1247 3262
rect 1281 3228 1314 3262
rect 1213 3172 1314 3228
rect 1213 3138 1247 3172
rect 1281 3138 1314 3172
rect 1213 3082 1314 3138
rect 1213 3048 1247 3082
rect 1281 3048 1314 3082
rect 1213 2992 1314 3048
rect 1213 2958 1247 2992
rect 1281 2958 1314 2992
rect 1213 2902 1314 2958
rect 1213 2868 1247 2902
rect 1281 2868 1314 2902
rect 1213 2812 1314 2868
rect 1213 2778 1247 2812
rect 1281 2778 1314 2812
rect 26 2688 60 2722
rect 94 2688 127 2722
rect 26 2673 127 2688
rect 1213 2722 1314 2778
rect 1213 2688 1247 2722
rect 1281 2688 1314 2722
rect 1213 2673 1314 2688
rect 26 2638 1314 2673
rect 26 2604 156 2638
rect 190 2604 246 2638
rect 280 2604 336 2638
rect 370 2604 426 2638
rect 460 2604 516 2638
rect 550 2604 606 2638
rect 640 2604 696 2638
rect 730 2604 786 2638
rect 820 2604 876 2638
rect 910 2604 966 2638
rect 1000 2604 1056 2638
rect 1090 2604 1146 2638
rect 1180 2604 1314 2638
rect 26 2572 1314 2604
rect 1368 3825 2656 3860
rect 1368 3802 1498 3825
rect 1368 3768 1402 3802
rect 1436 3791 1498 3802
rect 1532 3791 1588 3825
rect 1622 3791 1678 3825
rect 1712 3791 1768 3825
rect 1802 3791 1858 3825
rect 1892 3791 1948 3825
rect 1982 3791 2038 3825
rect 2072 3791 2128 3825
rect 2162 3791 2218 3825
rect 2252 3791 2308 3825
rect 2342 3791 2398 3825
rect 2432 3791 2488 3825
rect 2522 3802 2656 3825
rect 2522 3791 2589 3802
rect 1436 3768 2589 3791
rect 2623 3768 2656 3802
rect 1368 3759 2656 3768
rect 1368 3712 1469 3759
rect 1368 3678 1402 3712
rect 1436 3678 1469 3712
rect 2555 3712 2656 3759
rect 1368 3622 1469 3678
rect 1368 3588 1402 3622
rect 1436 3588 1469 3622
rect 1368 3532 1469 3588
rect 1368 3498 1402 3532
rect 1436 3498 1469 3532
rect 1368 3442 1469 3498
rect 1368 3408 1402 3442
rect 1436 3408 1469 3442
rect 1368 3352 1469 3408
rect 1368 3318 1402 3352
rect 1436 3318 1469 3352
rect 1368 3262 1469 3318
rect 1368 3228 1402 3262
rect 1436 3228 1469 3262
rect 1368 3172 1469 3228
rect 1368 3138 1402 3172
rect 1436 3138 1469 3172
rect 1368 3082 1469 3138
rect 1368 3048 1402 3082
rect 1436 3048 1469 3082
rect 1368 2992 1469 3048
rect 1368 2958 1402 2992
rect 1436 2958 1469 2992
rect 1368 2902 1469 2958
rect 1368 2868 1402 2902
rect 1436 2868 1469 2902
rect 1368 2812 1469 2868
rect 1368 2778 1402 2812
rect 1436 2778 1469 2812
rect 1368 2722 1469 2778
rect 2555 3678 2589 3712
rect 2623 3678 2656 3712
rect 2555 3622 2656 3678
rect 2555 3588 2589 3622
rect 2623 3588 2656 3622
rect 2555 3532 2656 3588
rect 2555 3498 2589 3532
rect 2623 3498 2656 3532
rect 2555 3442 2656 3498
rect 2555 3408 2589 3442
rect 2623 3408 2656 3442
rect 2555 3352 2656 3408
rect 2555 3318 2589 3352
rect 2623 3318 2656 3352
rect 2555 3262 2656 3318
rect 2555 3228 2589 3262
rect 2623 3228 2656 3262
rect 2555 3172 2656 3228
rect 2555 3138 2589 3172
rect 2623 3138 2656 3172
rect 2555 3082 2656 3138
rect 2555 3048 2589 3082
rect 2623 3048 2656 3082
rect 2555 2992 2656 3048
rect 2555 2958 2589 2992
rect 2623 2958 2656 2992
rect 2555 2902 2656 2958
rect 2555 2868 2589 2902
rect 2623 2868 2656 2902
rect 2555 2812 2656 2868
rect 2555 2778 2589 2812
rect 2623 2778 2656 2812
rect 1368 2688 1402 2722
rect 1436 2688 1469 2722
rect 1368 2673 1469 2688
rect 2555 2722 2656 2778
rect 2555 2688 2589 2722
rect 2623 2688 2656 2722
rect 2555 2673 2656 2688
rect 1368 2638 2656 2673
rect 1368 2604 1498 2638
rect 1532 2604 1588 2638
rect 1622 2604 1678 2638
rect 1712 2604 1768 2638
rect 1802 2604 1858 2638
rect 1892 2604 1948 2638
rect 1982 2604 2038 2638
rect 2072 2604 2128 2638
rect 2162 2604 2218 2638
rect 2252 2604 2308 2638
rect 2342 2604 2398 2638
rect 2432 2604 2488 2638
rect 2522 2604 2656 2638
rect 1368 2572 2656 2604
rect 2710 3825 3998 3860
rect 2710 3802 2840 3825
rect 2710 3768 2744 3802
rect 2778 3791 2840 3802
rect 2874 3791 2930 3825
rect 2964 3791 3020 3825
rect 3054 3791 3110 3825
rect 3144 3791 3200 3825
rect 3234 3791 3290 3825
rect 3324 3791 3380 3825
rect 3414 3791 3470 3825
rect 3504 3791 3560 3825
rect 3594 3791 3650 3825
rect 3684 3791 3740 3825
rect 3774 3791 3830 3825
rect 3864 3802 3998 3825
rect 3864 3791 3931 3802
rect 2778 3768 3931 3791
rect 3965 3768 3998 3802
rect 2710 3759 3998 3768
rect 2710 3712 2811 3759
rect 2710 3678 2744 3712
rect 2778 3678 2811 3712
rect 3897 3712 3998 3759
rect 2710 3622 2811 3678
rect 2710 3588 2744 3622
rect 2778 3588 2811 3622
rect 2710 3532 2811 3588
rect 2710 3498 2744 3532
rect 2778 3498 2811 3532
rect 2710 3442 2811 3498
rect 2710 3408 2744 3442
rect 2778 3408 2811 3442
rect 2710 3352 2811 3408
rect 2710 3318 2744 3352
rect 2778 3318 2811 3352
rect 2710 3262 2811 3318
rect 2710 3228 2744 3262
rect 2778 3228 2811 3262
rect 2710 3172 2811 3228
rect 2710 3138 2744 3172
rect 2778 3138 2811 3172
rect 2710 3082 2811 3138
rect 2710 3048 2744 3082
rect 2778 3048 2811 3082
rect 2710 2992 2811 3048
rect 2710 2958 2744 2992
rect 2778 2958 2811 2992
rect 2710 2902 2811 2958
rect 2710 2868 2744 2902
rect 2778 2868 2811 2902
rect 2710 2812 2811 2868
rect 2710 2778 2744 2812
rect 2778 2778 2811 2812
rect 2710 2722 2811 2778
rect 3897 3678 3931 3712
rect 3965 3678 3998 3712
rect 3897 3622 3998 3678
rect 3897 3588 3931 3622
rect 3965 3588 3998 3622
rect 3897 3532 3998 3588
rect 3897 3498 3931 3532
rect 3965 3498 3998 3532
rect 3897 3442 3998 3498
rect 3897 3408 3931 3442
rect 3965 3408 3998 3442
rect 3897 3352 3998 3408
rect 3897 3318 3931 3352
rect 3965 3318 3998 3352
rect 3897 3262 3998 3318
rect 3897 3228 3931 3262
rect 3965 3228 3998 3262
rect 3897 3172 3998 3228
rect 3897 3138 3931 3172
rect 3965 3138 3998 3172
rect 3897 3082 3998 3138
rect 3897 3048 3931 3082
rect 3965 3048 3998 3082
rect 3897 2992 3998 3048
rect 3897 2958 3931 2992
rect 3965 2958 3998 2992
rect 3897 2902 3998 2958
rect 3897 2868 3931 2902
rect 3965 2868 3998 2902
rect 3897 2812 3998 2868
rect 3897 2778 3931 2812
rect 3965 2778 3998 2812
rect 2710 2688 2744 2722
rect 2778 2688 2811 2722
rect 2710 2673 2811 2688
rect 3897 2722 3998 2778
rect 3897 2688 3931 2722
rect 3965 2688 3998 2722
rect 3897 2673 3998 2688
rect 2710 2638 3998 2673
rect 2710 2604 2840 2638
rect 2874 2604 2930 2638
rect 2964 2604 3020 2638
rect 3054 2604 3110 2638
rect 3144 2604 3200 2638
rect 3234 2604 3290 2638
rect 3324 2604 3380 2638
rect 3414 2604 3470 2638
rect 3504 2604 3560 2638
rect 3594 2604 3650 2638
rect 3684 2604 3740 2638
rect 3774 2604 3830 2638
rect 3864 2604 3998 2638
rect 2710 2572 3998 2604
rect 4052 3825 5340 3860
rect 4052 3802 4182 3825
rect 4052 3768 4086 3802
rect 4120 3791 4182 3802
rect 4216 3791 4272 3825
rect 4306 3791 4362 3825
rect 4396 3791 4452 3825
rect 4486 3791 4542 3825
rect 4576 3791 4632 3825
rect 4666 3791 4722 3825
rect 4756 3791 4812 3825
rect 4846 3791 4902 3825
rect 4936 3791 4992 3825
rect 5026 3791 5082 3825
rect 5116 3791 5172 3825
rect 5206 3802 5340 3825
rect 5206 3791 5273 3802
rect 4120 3768 5273 3791
rect 5307 3768 5340 3802
rect 4052 3759 5340 3768
rect 4052 3712 4153 3759
rect 4052 3678 4086 3712
rect 4120 3678 4153 3712
rect 5239 3712 5340 3759
rect 4052 3622 4153 3678
rect 4052 3588 4086 3622
rect 4120 3588 4153 3622
rect 4052 3532 4153 3588
rect 4052 3498 4086 3532
rect 4120 3498 4153 3532
rect 4052 3442 4153 3498
rect 4052 3408 4086 3442
rect 4120 3408 4153 3442
rect 4052 3352 4153 3408
rect 4052 3318 4086 3352
rect 4120 3318 4153 3352
rect 4052 3262 4153 3318
rect 4052 3228 4086 3262
rect 4120 3228 4153 3262
rect 4052 3172 4153 3228
rect 4052 3138 4086 3172
rect 4120 3138 4153 3172
rect 4052 3082 4153 3138
rect 4052 3048 4086 3082
rect 4120 3048 4153 3082
rect 4052 2992 4153 3048
rect 4052 2958 4086 2992
rect 4120 2958 4153 2992
rect 4052 2902 4153 2958
rect 4052 2868 4086 2902
rect 4120 2868 4153 2902
rect 4052 2812 4153 2868
rect 4052 2778 4086 2812
rect 4120 2778 4153 2812
rect 4052 2722 4153 2778
rect 5239 3678 5273 3712
rect 5307 3678 5340 3712
rect 5239 3622 5340 3678
rect 5239 3588 5273 3622
rect 5307 3588 5340 3622
rect 5239 3532 5340 3588
rect 5239 3498 5273 3532
rect 5307 3498 5340 3532
rect 5239 3442 5340 3498
rect 5239 3408 5273 3442
rect 5307 3408 5340 3442
rect 5239 3352 5340 3408
rect 5239 3318 5273 3352
rect 5307 3318 5340 3352
rect 5239 3262 5340 3318
rect 5239 3228 5273 3262
rect 5307 3228 5340 3262
rect 5239 3172 5340 3228
rect 5239 3138 5273 3172
rect 5307 3138 5340 3172
rect 5239 3082 5340 3138
rect 5239 3048 5273 3082
rect 5307 3048 5340 3082
rect 5239 2992 5340 3048
rect 5239 2958 5273 2992
rect 5307 2958 5340 2992
rect 5239 2902 5340 2958
rect 5239 2868 5273 2902
rect 5307 2868 5340 2902
rect 5239 2812 5340 2868
rect 5239 2778 5273 2812
rect 5307 2778 5340 2812
rect 4052 2688 4086 2722
rect 4120 2688 4153 2722
rect 4052 2673 4153 2688
rect 5239 2722 5340 2778
rect 5239 2688 5273 2722
rect 5307 2688 5340 2722
rect 5239 2673 5340 2688
rect 4052 2638 5340 2673
rect 4052 2604 4182 2638
rect 4216 2604 4272 2638
rect 4306 2604 4362 2638
rect 4396 2604 4452 2638
rect 4486 2604 4542 2638
rect 4576 2604 4632 2638
rect 4666 2604 4722 2638
rect 4756 2604 4812 2638
rect 4846 2604 4902 2638
rect 4936 2604 4992 2638
rect 5026 2604 5082 2638
rect 5116 2604 5172 2638
rect 5206 2604 5340 2638
rect 4052 2572 5340 2604
rect 5394 3825 6682 3860
rect 5394 3802 5524 3825
rect 5394 3768 5428 3802
rect 5462 3791 5524 3802
rect 5558 3791 5614 3825
rect 5648 3791 5704 3825
rect 5738 3791 5794 3825
rect 5828 3791 5884 3825
rect 5918 3791 5974 3825
rect 6008 3791 6064 3825
rect 6098 3791 6154 3825
rect 6188 3791 6244 3825
rect 6278 3791 6334 3825
rect 6368 3791 6424 3825
rect 6458 3791 6514 3825
rect 6548 3802 6682 3825
rect 6548 3791 6615 3802
rect 5462 3768 6615 3791
rect 6649 3768 6682 3802
rect 5394 3759 6682 3768
rect 5394 3712 5495 3759
rect 5394 3678 5428 3712
rect 5462 3678 5495 3712
rect 6581 3712 6682 3759
rect 5394 3622 5495 3678
rect 5394 3588 5428 3622
rect 5462 3588 5495 3622
rect 5394 3532 5495 3588
rect 5394 3498 5428 3532
rect 5462 3498 5495 3532
rect 5394 3442 5495 3498
rect 5394 3408 5428 3442
rect 5462 3408 5495 3442
rect 5394 3352 5495 3408
rect 5394 3318 5428 3352
rect 5462 3318 5495 3352
rect 5394 3262 5495 3318
rect 5394 3228 5428 3262
rect 5462 3228 5495 3262
rect 5394 3172 5495 3228
rect 5394 3138 5428 3172
rect 5462 3138 5495 3172
rect 5394 3082 5495 3138
rect 5394 3048 5428 3082
rect 5462 3048 5495 3082
rect 5394 2992 5495 3048
rect 5394 2958 5428 2992
rect 5462 2958 5495 2992
rect 5394 2902 5495 2958
rect 5394 2868 5428 2902
rect 5462 2868 5495 2902
rect 5394 2812 5495 2868
rect 5394 2778 5428 2812
rect 5462 2778 5495 2812
rect 5394 2722 5495 2778
rect 6581 3678 6615 3712
rect 6649 3678 6682 3712
rect 6581 3622 6682 3678
rect 6581 3588 6615 3622
rect 6649 3588 6682 3622
rect 6581 3532 6682 3588
rect 6581 3498 6615 3532
rect 6649 3498 6682 3532
rect 6581 3442 6682 3498
rect 6581 3408 6615 3442
rect 6649 3408 6682 3442
rect 6581 3352 6682 3408
rect 6581 3318 6615 3352
rect 6649 3318 6682 3352
rect 6581 3262 6682 3318
rect 6581 3228 6615 3262
rect 6649 3228 6682 3262
rect 6581 3172 6682 3228
rect 6581 3138 6615 3172
rect 6649 3138 6682 3172
rect 6581 3082 6682 3138
rect 6581 3048 6615 3082
rect 6649 3048 6682 3082
rect 6581 2992 6682 3048
rect 6581 2958 6615 2992
rect 6649 2958 6682 2992
rect 6581 2902 6682 2958
rect 6581 2868 6615 2902
rect 6649 2868 6682 2902
rect 6581 2812 6682 2868
rect 6581 2778 6615 2812
rect 6649 2778 6682 2812
rect 5394 2688 5428 2722
rect 5462 2688 5495 2722
rect 5394 2673 5495 2688
rect 6581 2722 6682 2778
rect 6581 2688 6615 2722
rect 6649 2688 6682 2722
rect 6581 2673 6682 2688
rect 5394 2638 6682 2673
rect 5394 2604 5524 2638
rect 5558 2604 5614 2638
rect 5648 2604 5704 2638
rect 5738 2604 5794 2638
rect 5828 2604 5884 2638
rect 5918 2604 5974 2638
rect 6008 2604 6064 2638
rect 6098 2604 6154 2638
rect 6188 2604 6244 2638
rect 6278 2604 6334 2638
rect 6368 2604 6424 2638
rect 6458 2604 6514 2638
rect 6548 2604 6682 2638
rect 5394 2572 6682 2604
rect 6736 3825 8024 3860
rect 6736 3802 6866 3825
rect 6736 3768 6770 3802
rect 6804 3791 6866 3802
rect 6900 3791 6956 3825
rect 6990 3791 7046 3825
rect 7080 3791 7136 3825
rect 7170 3791 7226 3825
rect 7260 3791 7316 3825
rect 7350 3791 7406 3825
rect 7440 3791 7496 3825
rect 7530 3791 7586 3825
rect 7620 3791 7676 3825
rect 7710 3791 7766 3825
rect 7800 3791 7856 3825
rect 7890 3802 8024 3825
rect 7890 3791 7957 3802
rect 6804 3768 7957 3791
rect 7991 3768 8024 3802
rect 6736 3759 8024 3768
rect 6736 3712 6837 3759
rect 6736 3678 6770 3712
rect 6804 3678 6837 3712
rect 7923 3712 8024 3759
rect 6736 3622 6837 3678
rect 6736 3588 6770 3622
rect 6804 3588 6837 3622
rect 6736 3532 6837 3588
rect 6736 3498 6770 3532
rect 6804 3498 6837 3532
rect 6736 3442 6837 3498
rect 6736 3408 6770 3442
rect 6804 3408 6837 3442
rect 6736 3352 6837 3408
rect 6736 3318 6770 3352
rect 6804 3318 6837 3352
rect 6736 3262 6837 3318
rect 6736 3228 6770 3262
rect 6804 3228 6837 3262
rect 6736 3172 6837 3228
rect 6736 3138 6770 3172
rect 6804 3138 6837 3172
rect 6736 3082 6837 3138
rect 6736 3048 6770 3082
rect 6804 3048 6837 3082
rect 6736 2992 6837 3048
rect 6736 2958 6770 2992
rect 6804 2958 6837 2992
rect 6736 2902 6837 2958
rect 6736 2868 6770 2902
rect 6804 2868 6837 2902
rect 6736 2812 6837 2868
rect 6736 2778 6770 2812
rect 6804 2778 6837 2812
rect 6736 2722 6837 2778
rect 7923 3678 7957 3712
rect 7991 3678 8024 3712
rect 7923 3622 8024 3678
rect 7923 3588 7957 3622
rect 7991 3588 8024 3622
rect 7923 3532 8024 3588
rect 7923 3498 7957 3532
rect 7991 3498 8024 3532
rect 7923 3442 8024 3498
rect 7923 3408 7957 3442
rect 7991 3408 8024 3442
rect 7923 3352 8024 3408
rect 7923 3318 7957 3352
rect 7991 3318 8024 3352
rect 7923 3262 8024 3318
rect 7923 3228 7957 3262
rect 7991 3228 8024 3262
rect 7923 3172 8024 3228
rect 7923 3138 7957 3172
rect 7991 3138 8024 3172
rect 7923 3082 8024 3138
rect 7923 3048 7957 3082
rect 7991 3048 8024 3082
rect 7923 2992 8024 3048
rect 7923 2958 7957 2992
rect 7991 2958 8024 2992
rect 7923 2902 8024 2958
rect 7923 2868 7957 2902
rect 7991 2868 8024 2902
rect 7923 2812 8024 2868
rect 7923 2778 7957 2812
rect 7991 2778 8024 2812
rect 6736 2688 6770 2722
rect 6804 2688 6837 2722
rect 6736 2673 6837 2688
rect 7923 2722 8024 2778
rect 7923 2688 7957 2722
rect 7991 2688 8024 2722
rect 7923 2673 8024 2688
rect 6736 2638 8024 2673
rect 6736 2604 6866 2638
rect 6900 2604 6956 2638
rect 6990 2604 7046 2638
rect 7080 2604 7136 2638
rect 7170 2604 7226 2638
rect 7260 2604 7316 2638
rect 7350 2604 7406 2638
rect 7440 2604 7496 2638
rect 7530 2604 7586 2638
rect 7620 2604 7676 2638
rect 7710 2604 7766 2638
rect 7800 2604 7856 2638
rect 7890 2604 8024 2638
rect 6736 2572 8024 2604
rect 8078 3825 9366 3860
rect 8078 3802 8208 3825
rect 8078 3768 8112 3802
rect 8146 3791 8208 3802
rect 8242 3791 8298 3825
rect 8332 3791 8388 3825
rect 8422 3791 8478 3825
rect 8512 3791 8568 3825
rect 8602 3791 8658 3825
rect 8692 3791 8748 3825
rect 8782 3791 8838 3825
rect 8872 3791 8928 3825
rect 8962 3791 9018 3825
rect 9052 3791 9108 3825
rect 9142 3791 9198 3825
rect 9232 3802 9366 3825
rect 9232 3791 9299 3802
rect 8146 3768 9299 3791
rect 9333 3768 9366 3802
rect 8078 3759 9366 3768
rect 8078 3712 8179 3759
rect 8078 3678 8112 3712
rect 8146 3678 8179 3712
rect 9265 3712 9366 3759
rect 8078 3622 8179 3678
rect 8078 3588 8112 3622
rect 8146 3588 8179 3622
rect 8078 3532 8179 3588
rect 8078 3498 8112 3532
rect 8146 3498 8179 3532
rect 8078 3442 8179 3498
rect 8078 3408 8112 3442
rect 8146 3408 8179 3442
rect 8078 3352 8179 3408
rect 8078 3318 8112 3352
rect 8146 3318 8179 3352
rect 8078 3262 8179 3318
rect 8078 3228 8112 3262
rect 8146 3228 8179 3262
rect 8078 3172 8179 3228
rect 8078 3138 8112 3172
rect 8146 3138 8179 3172
rect 8078 3082 8179 3138
rect 8078 3048 8112 3082
rect 8146 3048 8179 3082
rect 8078 2992 8179 3048
rect 8078 2958 8112 2992
rect 8146 2958 8179 2992
rect 8078 2902 8179 2958
rect 8078 2868 8112 2902
rect 8146 2868 8179 2902
rect 8078 2812 8179 2868
rect 8078 2778 8112 2812
rect 8146 2778 8179 2812
rect 8078 2722 8179 2778
rect 9265 3678 9299 3712
rect 9333 3678 9366 3712
rect 9265 3622 9366 3678
rect 9265 3588 9299 3622
rect 9333 3588 9366 3622
rect 9265 3532 9366 3588
rect 9265 3498 9299 3532
rect 9333 3498 9366 3532
rect 9265 3442 9366 3498
rect 9265 3408 9299 3442
rect 9333 3408 9366 3442
rect 9265 3352 9366 3408
rect 9265 3318 9299 3352
rect 9333 3318 9366 3352
rect 9265 3262 9366 3318
rect 9265 3228 9299 3262
rect 9333 3228 9366 3262
rect 9265 3172 9366 3228
rect 9265 3138 9299 3172
rect 9333 3138 9366 3172
rect 9265 3082 9366 3138
rect 9265 3048 9299 3082
rect 9333 3048 9366 3082
rect 9265 2992 9366 3048
rect 9265 2958 9299 2992
rect 9333 2958 9366 2992
rect 9265 2902 9366 2958
rect 9265 2868 9299 2902
rect 9333 2868 9366 2902
rect 9265 2812 9366 2868
rect 9265 2778 9299 2812
rect 9333 2778 9366 2812
rect 8078 2688 8112 2722
rect 8146 2688 8179 2722
rect 8078 2673 8179 2688
rect 9265 2722 9366 2778
rect 9265 2688 9299 2722
rect 9333 2688 9366 2722
rect 9265 2673 9366 2688
rect 8078 2638 9366 2673
rect 8078 2604 8208 2638
rect 8242 2604 8298 2638
rect 8332 2604 8388 2638
rect 8422 2604 8478 2638
rect 8512 2604 8568 2638
rect 8602 2604 8658 2638
rect 8692 2604 8748 2638
rect 8782 2604 8838 2638
rect 8872 2604 8928 2638
rect 8962 2604 9018 2638
rect 9052 2604 9108 2638
rect 9142 2604 9198 2638
rect 9232 2604 9366 2638
rect 8078 2572 9366 2604
rect 26 2483 1314 2518
rect 26 2460 156 2483
rect 26 2426 60 2460
rect 94 2449 156 2460
rect 190 2449 246 2483
rect 280 2449 336 2483
rect 370 2449 426 2483
rect 460 2449 516 2483
rect 550 2449 606 2483
rect 640 2449 696 2483
rect 730 2449 786 2483
rect 820 2449 876 2483
rect 910 2449 966 2483
rect 1000 2449 1056 2483
rect 1090 2449 1146 2483
rect 1180 2460 1314 2483
rect 1180 2449 1247 2460
rect 94 2426 1247 2449
rect 1281 2426 1314 2460
rect 26 2417 1314 2426
rect 26 2370 127 2417
rect 26 2336 60 2370
rect 94 2336 127 2370
rect 1213 2370 1314 2417
rect 26 2280 127 2336
rect 26 2246 60 2280
rect 94 2246 127 2280
rect 26 2190 127 2246
rect 26 2156 60 2190
rect 94 2156 127 2190
rect 26 2100 127 2156
rect 26 2066 60 2100
rect 94 2066 127 2100
rect 26 2010 127 2066
rect 26 1976 60 2010
rect 94 1976 127 2010
rect 26 1920 127 1976
rect 26 1886 60 1920
rect 94 1886 127 1920
rect 26 1830 127 1886
rect 26 1796 60 1830
rect 94 1796 127 1830
rect 26 1740 127 1796
rect 26 1706 60 1740
rect 94 1706 127 1740
rect 26 1650 127 1706
rect 26 1616 60 1650
rect 94 1616 127 1650
rect 26 1560 127 1616
rect 26 1526 60 1560
rect 94 1526 127 1560
rect 26 1470 127 1526
rect 26 1436 60 1470
rect 94 1436 127 1470
rect 26 1380 127 1436
rect 1213 2336 1247 2370
rect 1281 2336 1314 2370
rect 1213 2280 1314 2336
rect 1213 2246 1247 2280
rect 1281 2246 1314 2280
rect 1213 2190 1314 2246
rect 1213 2156 1247 2190
rect 1281 2156 1314 2190
rect 1213 2100 1314 2156
rect 1213 2066 1247 2100
rect 1281 2066 1314 2100
rect 1213 2010 1314 2066
rect 1213 1976 1247 2010
rect 1281 1976 1314 2010
rect 1213 1920 1314 1976
rect 1213 1886 1247 1920
rect 1281 1886 1314 1920
rect 1213 1830 1314 1886
rect 1213 1796 1247 1830
rect 1281 1796 1314 1830
rect 1213 1740 1314 1796
rect 1213 1706 1247 1740
rect 1281 1706 1314 1740
rect 1213 1650 1314 1706
rect 1213 1616 1247 1650
rect 1281 1616 1314 1650
rect 1213 1560 1314 1616
rect 1213 1526 1247 1560
rect 1281 1526 1314 1560
rect 1213 1470 1314 1526
rect 1213 1436 1247 1470
rect 1281 1436 1314 1470
rect 26 1346 60 1380
rect 94 1346 127 1380
rect 26 1331 127 1346
rect 1213 1380 1314 1436
rect 1213 1346 1247 1380
rect 1281 1346 1314 1380
rect 1213 1331 1314 1346
rect 26 1296 1314 1331
rect 26 1262 156 1296
rect 190 1262 246 1296
rect 280 1262 336 1296
rect 370 1262 426 1296
rect 460 1262 516 1296
rect 550 1262 606 1296
rect 640 1262 696 1296
rect 730 1262 786 1296
rect 820 1262 876 1296
rect 910 1262 966 1296
rect 1000 1262 1056 1296
rect 1090 1262 1146 1296
rect 1180 1262 1314 1296
rect 26 1230 1314 1262
rect 1368 2483 2656 2518
rect 1368 2460 1498 2483
rect 1368 2426 1402 2460
rect 1436 2449 1498 2460
rect 1532 2449 1588 2483
rect 1622 2449 1678 2483
rect 1712 2449 1768 2483
rect 1802 2449 1858 2483
rect 1892 2449 1948 2483
rect 1982 2449 2038 2483
rect 2072 2449 2128 2483
rect 2162 2449 2218 2483
rect 2252 2449 2308 2483
rect 2342 2449 2398 2483
rect 2432 2449 2488 2483
rect 2522 2460 2656 2483
rect 2522 2449 2589 2460
rect 1436 2426 2589 2449
rect 2623 2426 2656 2460
rect 1368 2417 2656 2426
rect 1368 2370 1469 2417
rect 1368 2336 1402 2370
rect 1436 2336 1469 2370
rect 2555 2370 2656 2417
rect 1368 2280 1469 2336
rect 1368 2246 1402 2280
rect 1436 2246 1469 2280
rect 1368 2190 1469 2246
rect 1368 2156 1402 2190
rect 1436 2156 1469 2190
rect 1368 2100 1469 2156
rect 1368 2066 1402 2100
rect 1436 2066 1469 2100
rect 1368 2010 1469 2066
rect 1368 1976 1402 2010
rect 1436 1976 1469 2010
rect 1368 1920 1469 1976
rect 1368 1886 1402 1920
rect 1436 1886 1469 1920
rect 1368 1830 1469 1886
rect 1368 1796 1402 1830
rect 1436 1796 1469 1830
rect 1368 1740 1469 1796
rect 1368 1706 1402 1740
rect 1436 1706 1469 1740
rect 1368 1650 1469 1706
rect 1368 1616 1402 1650
rect 1436 1616 1469 1650
rect 1368 1560 1469 1616
rect 1368 1526 1402 1560
rect 1436 1526 1469 1560
rect 1368 1470 1469 1526
rect 1368 1436 1402 1470
rect 1436 1436 1469 1470
rect 1368 1380 1469 1436
rect 2555 2336 2589 2370
rect 2623 2336 2656 2370
rect 2555 2280 2656 2336
rect 2555 2246 2589 2280
rect 2623 2246 2656 2280
rect 2555 2190 2656 2246
rect 2555 2156 2589 2190
rect 2623 2156 2656 2190
rect 2555 2100 2656 2156
rect 2555 2066 2589 2100
rect 2623 2066 2656 2100
rect 2555 2010 2656 2066
rect 2555 1976 2589 2010
rect 2623 1976 2656 2010
rect 2555 1920 2656 1976
rect 2555 1886 2589 1920
rect 2623 1886 2656 1920
rect 2555 1830 2656 1886
rect 2555 1796 2589 1830
rect 2623 1796 2656 1830
rect 2555 1740 2656 1796
rect 2555 1706 2589 1740
rect 2623 1706 2656 1740
rect 2555 1650 2656 1706
rect 2555 1616 2589 1650
rect 2623 1616 2656 1650
rect 2555 1560 2656 1616
rect 2555 1526 2589 1560
rect 2623 1526 2656 1560
rect 2555 1470 2656 1526
rect 2555 1436 2589 1470
rect 2623 1436 2656 1470
rect 1368 1346 1402 1380
rect 1436 1346 1469 1380
rect 1368 1331 1469 1346
rect 2555 1380 2656 1436
rect 2555 1346 2589 1380
rect 2623 1346 2656 1380
rect 2555 1331 2656 1346
rect 1368 1296 2656 1331
rect 1368 1262 1498 1296
rect 1532 1262 1588 1296
rect 1622 1262 1678 1296
rect 1712 1262 1768 1296
rect 1802 1262 1858 1296
rect 1892 1262 1948 1296
rect 1982 1262 2038 1296
rect 2072 1262 2128 1296
rect 2162 1262 2218 1296
rect 2252 1262 2308 1296
rect 2342 1262 2398 1296
rect 2432 1262 2488 1296
rect 2522 1262 2656 1296
rect 1368 1230 2656 1262
rect 2710 2483 3998 2518
rect 2710 2460 2840 2483
rect 2710 2426 2744 2460
rect 2778 2449 2840 2460
rect 2874 2449 2930 2483
rect 2964 2449 3020 2483
rect 3054 2449 3110 2483
rect 3144 2449 3200 2483
rect 3234 2449 3290 2483
rect 3324 2449 3380 2483
rect 3414 2449 3470 2483
rect 3504 2449 3560 2483
rect 3594 2449 3650 2483
rect 3684 2449 3740 2483
rect 3774 2449 3830 2483
rect 3864 2460 3998 2483
rect 3864 2449 3931 2460
rect 2778 2426 3931 2449
rect 3965 2426 3998 2460
rect 2710 2417 3998 2426
rect 2710 2370 2811 2417
rect 2710 2336 2744 2370
rect 2778 2336 2811 2370
rect 3897 2370 3998 2417
rect 2710 2280 2811 2336
rect 2710 2246 2744 2280
rect 2778 2246 2811 2280
rect 2710 2190 2811 2246
rect 2710 2156 2744 2190
rect 2778 2156 2811 2190
rect 2710 2100 2811 2156
rect 2710 2066 2744 2100
rect 2778 2066 2811 2100
rect 2710 2010 2811 2066
rect 2710 1976 2744 2010
rect 2778 1976 2811 2010
rect 2710 1920 2811 1976
rect 2710 1886 2744 1920
rect 2778 1886 2811 1920
rect 2710 1830 2811 1886
rect 2710 1796 2744 1830
rect 2778 1796 2811 1830
rect 2710 1740 2811 1796
rect 2710 1706 2744 1740
rect 2778 1706 2811 1740
rect 2710 1650 2811 1706
rect 2710 1616 2744 1650
rect 2778 1616 2811 1650
rect 2710 1560 2811 1616
rect 2710 1526 2744 1560
rect 2778 1526 2811 1560
rect 2710 1470 2811 1526
rect 2710 1436 2744 1470
rect 2778 1436 2811 1470
rect 2710 1380 2811 1436
rect 3897 2336 3931 2370
rect 3965 2336 3998 2370
rect 3897 2280 3998 2336
rect 3897 2246 3931 2280
rect 3965 2246 3998 2280
rect 3897 2190 3998 2246
rect 3897 2156 3931 2190
rect 3965 2156 3998 2190
rect 3897 2100 3998 2156
rect 3897 2066 3931 2100
rect 3965 2066 3998 2100
rect 3897 2010 3998 2066
rect 3897 1976 3931 2010
rect 3965 1976 3998 2010
rect 3897 1920 3998 1976
rect 3897 1886 3931 1920
rect 3965 1886 3998 1920
rect 3897 1830 3998 1886
rect 3897 1796 3931 1830
rect 3965 1796 3998 1830
rect 3897 1740 3998 1796
rect 3897 1706 3931 1740
rect 3965 1706 3998 1740
rect 3897 1650 3998 1706
rect 3897 1616 3931 1650
rect 3965 1616 3998 1650
rect 3897 1560 3998 1616
rect 3897 1526 3931 1560
rect 3965 1526 3998 1560
rect 3897 1470 3998 1526
rect 3897 1436 3931 1470
rect 3965 1436 3998 1470
rect 2710 1346 2744 1380
rect 2778 1346 2811 1380
rect 2710 1331 2811 1346
rect 3897 1380 3998 1436
rect 3897 1346 3931 1380
rect 3965 1346 3998 1380
rect 3897 1331 3998 1346
rect 2710 1296 3998 1331
rect 2710 1262 2840 1296
rect 2874 1262 2930 1296
rect 2964 1262 3020 1296
rect 3054 1262 3110 1296
rect 3144 1262 3200 1296
rect 3234 1262 3290 1296
rect 3324 1262 3380 1296
rect 3414 1262 3470 1296
rect 3504 1262 3560 1296
rect 3594 1262 3650 1296
rect 3684 1262 3740 1296
rect 3774 1262 3830 1296
rect 3864 1262 3998 1296
rect 2710 1230 3998 1262
rect 4052 2483 5340 2518
rect 4052 2460 4182 2483
rect 4052 2426 4086 2460
rect 4120 2449 4182 2460
rect 4216 2449 4272 2483
rect 4306 2449 4362 2483
rect 4396 2449 4452 2483
rect 4486 2449 4542 2483
rect 4576 2449 4632 2483
rect 4666 2449 4722 2483
rect 4756 2449 4812 2483
rect 4846 2449 4902 2483
rect 4936 2449 4992 2483
rect 5026 2449 5082 2483
rect 5116 2449 5172 2483
rect 5206 2460 5340 2483
rect 5206 2449 5273 2460
rect 4120 2426 5273 2449
rect 5307 2426 5340 2460
rect 4052 2417 5340 2426
rect 4052 2370 4153 2417
rect 4052 2336 4086 2370
rect 4120 2336 4153 2370
rect 5239 2370 5340 2417
rect 4052 2280 4153 2336
rect 4052 2246 4086 2280
rect 4120 2246 4153 2280
rect 4052 2190 4153 2246
rect 4052 2156 4086 2190
rect 4120 2156 4153 2190
rect 4052 2100 4153 2156
rect 4052 2066 4086 2100
rect 4120 2066 4153 2100
rect 4052 2010 4153 2066
rect 4052 1976 4086 2010
rect 4120 1976 4153 2010
rect 4052 1920 4153 1976
rect 4052 1886 4086 1920
rect 4120 1886 4153 1920
rect 4052 1830 4153 1886
rect 4052 1796 4086 1830
rect 4120 1796 4153 1830
rect 4052 1740 4153 1796
rect 4052 1706 4086 1740
rect 4120 1706 4153 1740
rect 4052 1650 4153 1706
rect 4052 1616 4086 1650
rect 4120 1616 4153 1650
rect 4052 1560 4153 1616
rect 4052 1526 4086 1560
rect 4120 1526 4153 1560
rect 4052 1470 4153 1526
rect 4052 1436 4086 1470
rect 4120 1436 4153 1470
rect 4052 1380 4153 1436
rect 5239 2336 5273 2370
rect 5307 2336 5340 2370
rect 5239 2280 5340 2336
rect 5239 2246 5273 2280
rect 5307 2246 5340 2280
rect 5239 2190 5340 2246
rect 5239 2156 5273 2190
rect 5307 2156 5340 2190
rect 5239 2100 5340 2156
rect 5239 2066 5273 2100
rect 5307 2066 5340 2100
rect 5239 2010 5340 2066
rect 5239 1976 5273 2010
rect 5307 1976 5340 2010
rect 5239 1920 5340 1976
rect 5239 1886 5273 1920
rect 5307 1886 5340 1920
rect 5239 1830 5340 1886
rect 5239 1796 5273 1830
rect 5307 1796 5340 1830
rect 5239 1740 5340 1796
rect 5239 1706 5273 1740
rect 5307 1706 5340 1740
rect 5239 1650 5340 1706
rect 5239 1616 5273 1650
rect 5307 1616 5340 1650
rect 5239 1560 5340 1616
rect 5239 1526 5273 1560
rect 5307 1526 5340 1560
rect 5239 1470 5340 1526
rect 5239 1436 5273 1470
rect 5307 1436 5340 1470
rect 4052 1346 4086 1380
rect 4120 1346 4153 1380
rect 4052 1331 4153 1346
rect 5239 1380 5340 1436
rect 5239 1346 5273 1380
rect 5307 1346 5340 1380
rect 5239 1331 5340 1346
rect 4052 1296 5340 1331
rect 4052 1262 4182 1296
rect 4216 1262 4272 1296
rect 4306 1262 4362 1296
rect 4396 1262 4452 1296
rect 4486 1262 4542 1296
rect 4576 1262 4632 1296
rect 4666 1262 4722 1296
rect 4756 1262 4812 1296
rect 4846 1262 4902 1296
rect 4936 1262 4992 1296
rect 5026 1262 5082 1296
rect 5116 1262 5172 1296
rect 5206 1262 5340 1296
rect 4052 1230 5340 1262
rect 5394 2483 6682 2518
rect 5394 2460 5524 2483
rect 5394 2426 5428 2460
rect 5462 2449 5524 2460
rect 5558 2449 5614 2483
rect 5648 2449 5704 2483
rect 5738 2449 5794 2483
rect 5828 2449 5884 2483
rect 5918 2449 5974 2483
rect 6008 2449 6064 2483
rect 6098 2449 6154 2483
rect 6188 2449 6244 2483
rect 6278 2449 6334 2483
rect 6368 2449 6424 2483
rect 6458 2449 6514 2483
rect 6548 2460 6682 2483
rect 6548 2449 6615 2460
rect 5462 2426 6615 2449
rect 6649 2426 6682 2460
rect 5394 2417 6682 2426
rect 5394 2370 5495 2417
rect 5394 2336 5428 2370
rect 5462 2336 5495 2370
rect 6581 2370 6682 2417
rect 5394 2280 5495 2336
rect 5394 2246 5428 2280
rect 5462 2246 5495 2280
rect 5394 2190 5495 2246
rect 5394 2156 5428 2190
rect 5462 2156 5495 2190
rect 5394 2100 5495 2156
rect 5394 2066 5428 2100
rect 5462 2066 5495 2100
rect 5394 2010 5495 2066
rect 5394 1976 5428 2010
rect 5462 1976 5495 2010
rect 5394 1920 5495 1976
rect 5394 1886 5428 1920
rect 5462 1886 5495 1920
rect 5394 1830 5495 1886
rect 5394 1796 5428 1830
rect 5462 1796 5495 1830
rect 5394 1740 5495 1796
rect 5394 1706 5428 1740
rect 5462 1706 5495 1740
rect 5394 1650 5495 1706
rect 5394 1616 5428 1650
rect 5462 1616 5495 1650
rect 5394 1560 5495 1616
rect 5394 1526 5428 1560
rect 5462 1526 5495 1560
rect 5394 1470 5495 1526
rect 5394 1436 5428 1470
rect 5462 1436 5495 1470
rect 5394 1380 5495 1436
rect 6581 2336 6615 2370
rect 6649 2336 6682 2370
rect 6581 2280 6682 2336
rect 6581 2246 6615 2280
rect 6649 2246 6682 2280
rect 6581 2190 6682 2246
rect 6581 2156 6615 2190
rect 6649 2156 6682 2190
rect 6581 2100 6682 2156
rect 6581 2066 6615 2100
rect 6649 2066 6682 2100
rect 6581 2010 6682 2066
rect 6581 1976 6615 2010
rect 6649 1976 6682 2010
rect 6581 1920 6682 1976
rect 6581 1886 6615 1920
rect 6649 1886 6682 1920
rect 6581 1830 6682 1886
rect 6581 1796 6615 1830
rect 6649 1796 6682 1830
rect 6581 1740 6682 1796
rect 6581 1706 6615 1740
rect 6649 1706 6682 1740
rect 6581 1650 6682 1706
rect 6581 1616 6615 1650
rect 6649 1616 6682 1650
rect 6581 1560 6682 1616
rect 6581 1526 6615 1560
rect 6649 1526 6682 1560
rect 6581 1470 6682 1526
rect 6581 1436 6615 1470
rect 6649 1436 6682 1470
rect 5394 1346 5428 1380
rect 5462 1346 5495 1380
rect 5394 1331 5495 1346
rect 6581 1380 6682 1436
rect 6581 1346 6615 1380
rect 6649 1346 6682 1380
rect 6581 1331 6682 1346
rect 5394 1296 6682 1331
rect 5394 1262 5524 1296
rect 5558 1262 5614 1296
rect 5648 1262 5704 1296
rect 5738 1262 5794 1296
rect 5828 1262 5884 1296
rect 5918 1262 5974 1296
rect 6008 1262 6064 1296
rect 6098 1262 6154 1296
rect 6188 1262 6244 1296
rect 6278 1262 6334 1296
rect 6368 1262 6424 1296
rect 6458 1262 6514 1296
rect 6548 1262 6682 1296
rect 5394 1230 6682 1262
rect 6736 2483 8024 2518
rect 6736 2460 6866 2483
rect 6736 2426 6770 2460
rect 6804 2449 6866 2460
rect 6900 2449 6956 2483
rect 6990 2449 7046 2483
rect 7080 2449 7136 2483
rect 7170 2449 7226 2483
rect 7260 2449 7316 2483
rect 7350 2449 7406 2483
rect 7440 2449 7496 2483
rect 7530 2449 7586 2483
rect 7620 2449 7676 2483
rect 7710 2449 7766 2483
rect 7800 2449 7856 2483
rect 7890 2460 8024 2483
rect 7890 2449 7957 2460
rect 6804 2426 7957 2449
rect 7991 2426 8024 2460
rect 6736 2417 8024 2426
rect 6736 2370 6837 2417
rect 6736 2336 6770 2370
rect 6804 2336 6837 2370
rect 7923 2370 8024 2417
rect 6736 2280 6837 2336
rect 6736 2246 6770 2280
rect 6804 2246 6837 2280
rect 6736 2190 6837 2246
rect 6736 2156 6770 2190
rect 6804 2156 6837 2190
rect 6736 2100 6837 2156
rect 6736 2066 6770 2100
rect 6804 2066 6837 2100
rect 6736 2010 6837 2066
rect 6736 1976 6770 2010
rect 6804 1976 6837 2010
rect 6736 1920 6837 1976
rect 6736 1886 6770 1920
rect 6804 1886 6837 1920
rect 6736 1830 6837 1886
rect 6736 1796 6770 1830
rect 6804 1796 6837 1830
rect 6736 1740 6837 1796
rect 6736 1706 6770 1740
rect 6804 1706 6837 1740
rect 6736 1650 6837 1706
rect 6736 1616 6770 1650
rect 6804 1616 6837 1650
rect 6736 1560 6837 1616
rect 6736 1526 6770 1560
rect 6804 1526 6837 1560
rect 6736 1470 6837 1526
rect 6736 1436 6770 1470
rect 6804 1436 6837 1470
rect 6736 1380 6837 1436
rect 7923 2336 7957 2370
rect 7991 2336 8024 2370
rect 7923 2280 8024 2336
rect 7923 2246 7957 2280
rect 7991 2246 8024 2280
rect 7923 2190 8024 2246
rect 7923 2156 7957 2190
rect 7991 2156 8024 2190
rect 7923 2100 8024 2156
rect 7923 2066 7957 2100
rect 7991 2066 8024 2100
rect 7923 2010 8024 2066
rect 7923 1976 7957 2010
rect 7991 1976 8024 2010
rect 7923 1920 8024 1976
rect 7923 1886 7957 1920
rect 7991 1886 8024 1920
rect 7923 1830 8024 1886
rect 7923 1796 7957 1830
rect 7991 1796 8024 1830
rect 7923 1740 8024 1796
rect 7923 1706 7957 1740
rect 7991 1706 8024 1740
rect 7923 1650 8024 1706
rect 7923 1616 7957 1650
rect 7991 1616 8024 1650
rect 7923 1560 8024 1616
rect 7923 1526 7957 1560
rect 7991 1526 8024 1560
rect 7923 1470 8024 1526
rect 7923 1436 7957 1470
rect 7991 1436 8024 1470
rect 6736 1346 6770 1380
rect 6804 1346 6837 1380
rect 6736 1331 6837 1346
rect 7923 1380 8024 1436
rect 7923 1346 7957 1380
rect 7991 1346 8024 1380
rect 7923 1331 8024 1346
rect 6736 1296 8024 1331
rect 6736 1262 6866 1296
rect 6900 1262 6956 1296
rect 6990 1262 7046 1296
rect 7080 1262 7136 1296
rect 7170 1262 7226 1296
rect 7260 1262 7316 1296
rect 7350 1262 7406 1296
rect 7440 1262 7496 1296
rect 7530 1262 7586 1296
rect 7620 1262 7676 1296
rect 7710 1262 7766 1296
rect 7800 1262 7856 1296
rect 7890 1262 8024 1296
rect 6736 1230 8024 1262
rect 8078 2483 9366 2518
rect 8078 2460 8208 2483
rect 8078 2426 8112 2460
rect 8146 2449 8208 2460
rect 8242 2449 8298 2483
rect 8332 2449 8388 2483
rect 8422 2449 8478 2483
rect 8512 2449 8568 2483
rect 8602 2449 8658 2483
rect 8692 2449 8748 2483
rect 8782 2449 8838 2483
rect 8872 2449 8928 2483
rect 8962 2449 9018 2483
rect 9052 2449 9108 2483
rect 9142 2449 9198 2483
rect 9232 2460 9366 2483
rect 9232 2449 9299 2460
rect 8146 2426 9299 2449
rect 9333 2426 9366 2460
rect 8078 2417 9366 2426
rect 8078 2370 8179 2417
rect 8078 2336 8112 2370
rect 8146 2336 8179 2370
rect 9265 2370 9366 2417
rect 8078 2280 8179 2336
rect 8078 2246 8112 2280
rect 8146 2246 8179 2280
rect 8078 2190 8179 2246
rect 8078 2156 8112 2190
rect 8146 2156 8179 2190
rect 8078 2100 8179 2156
rect 8078 2066 8112 2100
rect 8146 2066 8179 2100
rect 8078 2010 8179 2066
rect 8078 1976 8112 2010
rect 8146 1976 8179 2010
rect 8078 1920 8179 1976
rect 8078 1886 8112 1920
rect 8146 1886 8179 1920
rect 8078 1830 8179 1886
rect 8078 1796 8112 1830
rect 8146 1796 8179 1830
rect 8078 1740 8179 1796
rect 8078 1706 8112 1740
rect 8146 1706 8179 1740
rect 8078 1650 8179 1706
rect 8078 1616 8112 1650
rect 8146 1616 8179 1650
rect 8078 1560 8179 1616
rect 8078 1526 8112 1560
rect 8146 1526 8179 1560
rect 8078 1470 8179 1526
rect 8078 1436 8112 1470
rect 8146 1436 8179 1470
rect 8078 1380 8179 1436
rect 9265 2336 9299 2370
rect 9333 2336 9366 2370
rect 9265 2280 9366 2336
rect 9265 2246 9299 2280
rect 9333 2246 9366 2280
rect 9265 2190 9366 2246
rect 9265 2156 9299 2190
rect 9333 2156 9366 2190
rect 9265 2100 9366 2156
rect 9265 2066 9299 2100
rect 9333 2066 9366 2100
rect 9265 2010 9366 2066
rect 9265 1976 9299 2010
rect 9333 1976 9366 2010
rect 9265 1920 9366 1976
rect 9265 1886 9299 1920
rect 9333 1886 9366 1920
rect 9265 1830 9366 1886
rect 9265 1796 9299 1830
rect 9333 1796 9366 1830
rect 9265 1740 9366 1796
rect 9265 1706 9299 1740
rect 9333 1706 9366 1740
rect 9265 1650 9366 1706
rect 9265 1616 9299 1650
rect 9333 1616 9366 1650
rect 9265 1560 9366 1616
rect 9265 1526 9299 1560
rect 9333 1526 9366 1560
rect 9265 1470 9366 1526
rect 9265 1436 9299 1470
rect 9333 1436 9366 1470
rect 8078 1346 8112 1380
rect 8146 1346 8179 1380
rect 8078 1331 8179 1346
rect 9265 1380 9366 1436
rect 9265 1346 9299 1380
rect 9333 1346 9366 1380
rect 9265 1331 9366 1346
rect 8078 1296 9366 1331
rect 8078 1262 8208 1296
rect 8242 1262 8298 1296
rect 8332 1262 8388 1296
rect 8422 1262 8478 1296
rect 8512 1262 8568 1296
rect 8602 1262 8658 1296
rect 8692 1262 8748 1296
rect 8782 1262 8838 1296
rect 8872 1262 8928 1296
rect 8962 1262 9018 1296
rect 9052 1262 9108 1296
rect 9142 1262 9198 1296
rect 9232 1262 9366 1296
rect 8078 1230 9366 1262
rect 1686 1075 2656 1176
rect 1368 -11 1469 874
rect 2555 -11 2656 1075
rect 1368 -112 2656 -11
rect 2710 1075 3998 1176
rect 2710 -11 2811 1075
rect 3897 -11 3998 1075
rect 2710 -112 3998 -11
rect 4052 1075 5340 1176
rect 4052 -11 4153 1075
rect 5239 -11 5340 1075
rect 4052 -112 5340 -11
rect 5394 1075 6682 1176
rect 5394 -11 5495 1075
rect 6581 -11 6682 1075
rect 5394 -112 6682 -11
rect 6736 1141 8024 1176
rect 6736 1118 6866 1141
rect 6736 1084 6770 1118
rect 6804 1107 6866 1118
rect 6900 1107 6956 1141
rect 6990 1107 7046 1141
rect 7080 1107 7136 1141
rect 7170 1107 7226 1141
rect 7260 1107 7316 1141
rect 7350 1107 7406 1141
rect 7440 1107 7496 1141
rect 7530 1107 7586 1141
rect 7620 1107 7676 1141
rect 7710 1107 7766 1141
rect 7800 1107 7856 1141
rect 7890 1118 8024 1141
rect 7890 1107 7957 1118
rect 6804 1084 7957 1107
rect 7991 1084 8024 1118
rect 6736 1075 8024 1084
rect 6736 1028 6837 1075
rect 6736 994 6770 1028
rect 6804 994 6837 1028
rect 7923 1028 8024 1075
rect 6736 938 6837 994
rect 6736 904 6770 938
rect 6804 904 6837 938
rect 6736 848 6837 904
rect 6736 814 6770 848
rect 6804 814 6837 848
rect 6736 758 6837 814
rect 6736 724 6770 758
rect 6804 724 6837 758
rect 6736 668 6837 724
rect 6736 634 6770 668
rect 6804 634 6837 668
rect 6736 578 6837 634
rect 6736 544 6770 578
rect 6804 544 6837 578
rect 6736 488 6837 544
rect 6736 454 6770 488
rect 6804 454 6837 488
rect 6736 398 6837 454
rect 6736 364 6770 398
rect 6804 364 6837 398
rect 6736 308 6837 364
rect 6736 274 6770 308
rect 6804 274 6837 308
rect 6736 218 6837 274
rect 6736 184 6770 218
rect 6804 184 6837 218
rect 6736 128 6837 184
rect 6736 94 6770 128
rect 6804 94 6837 128
rect 6736 38 6837 94
rect 7923 994 7957 1028
rect 7991 994 8024 1028
rect 7923 938 8024 994
rect 7923 904 7957 938
rect 7991 904 8024 938
rect 7923 848 8024 904
rect 7923 814 7957 848
rect 7991 814 8024 848
rect 7923 758 8024 814
rect 7923 724 7957 758
rect 7991 724 8024 758
rect 7923 668 8024 724
rect 7923 634 7957 668
rect 7991 634 8024 668
rect 7923 578 8024 634
rect 7923 544 7957 578
rect 7991 544 8024 578
rect 7923 488 8024 544
rect 7923 454 7957 488
rect 7991 454 8024 488
rect 7923 398 8024 454
rect 7923 364 7957 398
rect 7991 364 8024 398
rect 7923 308 8024 364
rect 7923 274 7957 308
rect 7991 274 8024 308
rect 7923 218 8024 274
rect 7923 184 7957 218
rect 7991 184 8024 218
rect 7923 128 8024 184
rect 7923 94 7957 128
rect 7991 94 8024 128
rect 6736 4 6770 38
rect 6804 4 6837 38
rect 6736 -11 6837 4
rect 7923 38 8024 94
rect 7923 4 7957 38
rect 7991 4 8024 38
rect 7923 -11 8024 4
rect 6736 -46 8024 -11
rect 6736 -80 6866 -46
rect 6900 -80 6956 -46
rect 6990 -80 7046 -46
rect 7080 -80 7136 -46
rect 7170 -80 7226 -46
rect 7260 -80 7316 -46
rect 7350 -80 7406 -46
rect 7440 -80 7496 -46
rect 7530 -80 7586 -46
rect 7620 -80 7676 -46
rect 7710 -80 7766 -46
rect 7800 -80 7856 -46
rect 7890 -80 8024 -46
rect 6736 -112 8024 -80
rect 8078 1141 9366 1176
rect 8078 1118 8208 1141
rect 8078 1084 8112 1118
rect 8146 1107 8208 1118
rect 8242 1107 8298 1141
rect 8332 1107 8388 1141
rect 8422 1107 8478 1141
rect 8512 1107 8568 1141
rect 8602 1107 8658 1141
rect 8692 1107 8748 1141
rect 8782 1107 8838 1141
rect 8872 1107 8928 1141
rect 8962 1107 9018 1141
rect 9052 1107 9108 1141
rect 9142 1107 9198 1141
rect 9232 1118 9366 1141
rect 9232 1107 9299 1118
rect 8146 1084 9299 1107
rect 9333 1084 9366 1118
rect 8078 1075 9366 1084
rect 8078 1028 8179 1075
rect 8078 994 8112 1028
rect 8146 994 8179 1028
rect 9265 1028 9366 1075
rect 8078 938 8179 994
rect 8078 904 8112 938
rect 8146 904 8179 938
rect 8078 848 8179 904
rect 8078 814 8112 848
rect 8146 814 8179 848
rect 8078 758 8179 814
rect 8078 724 8112 758
rect 8146 724 8179 758
rect 8078 668 8179 724
rect 8078 634 8112 668
rect 8146 634 8179 668
rect 8078 578 8179 634
rect 8078 544 8112 578
rect 8146 544 8179 578
rect 8078 488 8179 544
rect 8078 454 8112 488
rect 8146 454 8179 488
rect 8078 398 8179 454
rect 8078 364 8112 398
rect 8146 364 8179 398
rect 8078 308 8179 364
rect 8078 274 8112 308
rect 8146 274 8179 308
rect 8078 218 8179 274
rect 8078 184 8112 218
rect 8146 184 8179 218
rect 8078 128 8179 184
rect 8078 94 8112 128
rect 8146 94 8179 128
rect 8078 38 8179 94
rect 9265 994 9299 1028
rect 9333 994 9366 1028
rect 9265 938 9366 994
rect 9265 904 9299 938
rect 9333 904 9366 938
rect 9265 848 9366 904
rect 9265 814 9299 848
rect 9333 814 9366 848
rect 9265 758 9366 814
rect 9265 724 9299 758
rect 9333 724 9366 758
rect 9265 668 9366 724
rect 9265 634 9299 668
rect 9333 634 9366 668
rect 9265 578 9366 634
rect 9265 544 9299 578
rect 9333 544 9366 578
rect 9265 488 9366 544
rect 9265 454 9299 488
rect 9333 454 9366 488
rect 9265 398 9366 454
rect 9265 364 9299 398
rect 9333 364 9366 398
rect 9265 308 9366 364
rect 9265 274 9299 308
rect 9333 274 9366 308
rect 9265 218 9366 274
rect 9265 184 9299 218
rect 9333 184 9366 218
rect 9265 128 9366 184
rect 9265 94 9299 128
rect 9333 94 9366 128
rect 8078 4 8112 38
rect 8146 4 8179 38
rect 8078 -11 8179 4
rect 9265 38 9366 94
rect 9265 4 9299 38
rect 9333 4 9366 38
rect 9265 -11 9366 4
rect 8078 -46 9366 -11
rect 8078 -80 8208 -46
rect 8242 -80 8298 -46
rect 8332 -80 8388 -46
rect 8422 -80 8478 -46
rect 8512 -80 8568 -46
rect 8602 -80 8658 -46
rect 8692 -80 8748 -46
rect 8782 -80 8838 -46
rect 8872 -80 8928 -46
rect 8962 -80 9018 -46
rect 9052 -80 9108 -46
rect 9142 -80 9198 -46
rect 9232 -80 9366 -46
rect 8078 -112 9366 -80
rect 26 -267 1314 -166
rect 26 -1353 127 -267
rect 1213 -1353 1314 -267
rect 26 -1454 1314 -1353
rect 1368 -267 2656 -166
rect 1368 -1353 1469 -267
rect 2555 -1353 2656 -267
rect 1368 -1454 2656 -1353
rect 2710 -267 3998 -166
rect 2710 -1353 2811 -267
rect 3897 -1353 3998 -267
rect 2710 -1454 3998 -1353
rect 4052 -267 5340 -166
rect 4052 -1353 4153 -267
rect 5239 -1353 5340 -267
rect 4052 -1454 5340 -1353
rect 5394 -267 6682 -166
rect 5394 -1353 5495 -267
rect 6581 -1353 6682 -267
rect 5394 -1454 6682 -1353
rect 6736 -201 8024 -166
rect 6736 -224 6866 -201
rect 6736 -258 6770 -224
rect 6804 -235 6866 -224
rect 6900 -235 6956 -201
rect 6990 -235 7046 -201
rect 7080 -235 7136 -201
rect 7170 -235 7226 -201
rect 7260 -235 7316 -201
rect 7350 -235 7406 -201
rect 7440 -235 7496 -201
rect 7530 -235 7586 -201
rect 7620 -235 7676 -201
rect 7710 -235 7766 -201
rect 7800 -235 7856 -201
rect 7890 -224 8024 -201
rect 7890 -235 7957 -224
rect 6804 -258 7957 -235
rect 7991 -258 8024 -224
rect 6736 -267 8024 -258
rect 6736 -314 6837 -267
rect 6736 -348 6770 -314
rect 6804 -348 6837 -314
rect 7923 -314 8024 -267
rect 6736 -404 6837 -348
rect 6736 -438 6770 -404
rect 6804 -438 6837 -404
rect 6736 -494 6837 -438
rect 6736 -528 6770 -494
rect 6804 -528 6837 -494
rect 6736 -584 6837 -528
rect 6736 -618 6770 -584
rect 6804 -618 6837 -584
rect 6736 -674 6837 -618
rect 6736 -708 6770 -674
rect 6804 -708 6837 -674
rect 6736 -764 6837 -708
rect 6736 -798 6770 -764
rect 6804 -798 6837 -764
rect 6736 -854 6837 -798
rect 6736 -888 6770 -854
rect 6804 -888 6837 -854
rect 6736 -944 6837 -888
rect 6736 -978 6770 -944
rect 6804 -978 6837 -944
rect 6736 -1034 6837 -978
rect 6736 -1068 6770 -1034
rect 6804 -1068 6837 -1034
rect 6736 -1124 6837 -1068
rect 6736 -1158 6770 -1124
rect 6804 -1158 6837 -1124
rect 6736 -1214 6837 -1158
rect 6736 -1248 6770 -1214
rect 6804 -1248 6837 -1214
rect 6736 -1304 6837 -1248
rect 7923 -348 7957 -314
rect 7991 -348 8024 -314
rect 7923 -404 8024 -348
rect 7923 -438 7957 -404
rect 7991 -438 8024 -404
rect 7923 -494 8024 -438
rect 7923 -528 7957 -494
rect 7991 -528 8024 -494
rect 7923 -584 8024 -528
rect 7923 -618 7957 -584
rect 7991 -618 8024 -584
rect 7923 -674 8024 -618
rect 7923 -708 7957 -674
rect 7991 -708 8024 -674
rect 7923 -764 8024 -708
rect 7923 -798 7957 -764
rect 7991 -798 8024 -764
rect 7923 -854 8024 -798
rect 7923 -888 7957 -854
rect 7991 -888 8024 -854
rect 7923 -944 8024 -888
rect 7923 -978 7957 -944
rect 7991 -978 8024 -944
rect 7923 -1034 8024 -978
rect 7923 -1068 7957 -1034
rect 7991 -1068 8024 -1034
rect 7923 -1124 8024 -1068
rect 7923 -1158 7957 -1124
rect 7991 -1158 8024 -1124
rect 7923 -1214 8024 -1158
rect 7923 -1248 7957 -1214
rect 7991 -1248 8024 -1214
rect 6736 -1338 6770 -1304
rect 6804 -1338 6837 -1304
rect 6736 -1353 6837 -1338
rect 7923 -1304 8024 -1248
rect 7923 -1338 7957 -1304
rect 7991 -1338 8024 -1304
rect 7923 -1353 8024 -1338
rect 6736 -1388 8024 -1353
rect 6736 -1422 6866 -1388
rect 6900 -1422 6956 -1388
rect 6990 -1422 7046 -1388
rect 7080 -1422 7136 -1388
rect 7170 -1422 7226 -1388
rect 7260 -1422 7316 -1388
rect 7350 -1422 7406 -1388
rect 7440 -1422 7496 -1388
rect 7530 -1422 7586 -1388
rect 7620 -1422 7676 -1388
rect 7710 -1422 7766 -1388
rect 7800 -1422 7856 -1388
rect 7890 -1422 8024 -1388
rect 6736 -1454 8024 -1422
rect 8078 -201 9366 -166
rect 8078 -224 8208 -201
rect 8078 -258 8112 -224
rect 8146 -235 8208 -224
rect 8242 -235 8298 -201
rect 8332 -235 8388 -201
rect 8422 -235 8478 -201
rect 8512 -235 8568 -201
rect 8602 -235 8658 -201
rect 8692 -235 8748 -201
rect 8782 -235 8838 -201
rect 8872 -235 8928 -201
rect 8962 -235 9018 -201
rect 9052 -235 9108 -201
rect 9142 -235 9198 -201
rect 9232 -224 9366 -201
rect 9232 -235 9299 -224
rect 8146 -258 9299 -235
rect 9333 -258 9366 -224
rect 8078 -267 9366 -258
rect 8078 -314 8179 -267
rect 8078 -348 8112 -314
rect 8146 -348 8179 -314
rect 9265 -314 9366 -267
rect 8078 -404 8179 -348
rect 8078 -438 8112 -404
rect 8146 -438 8179 -404
rect 8078 -494 8179 -438
rect 8078 -528 8112 -494
rect 8146 -528 8179 -494
rect 8078 -584 8179 -528
rect 8078 -618 8112 -584
rect 8146 -618 8179 -584
rect 8078 -674 8179 -618
rect 8078 -708 8112 -674
rect 8146 -708 8179 -674
rect 8078 -764 8179 -708
rect 8078 -798 8112 -764
rect 8146 -798 8179 -764
rect 8078 -854 8179 -798
rect 8078 -888 8112 -854
rect 8146 -888 8179 -854
rect 8078 -944 8179 -888
rect 8078 -978 8112 -944
rect 8146 -978 8179 -944
rect 8078 -1034 8179 -978
rect 8078 -1068 8112 -1034
rect 8146 -1068 8179 -1034
rect 8078 -1124 8179 -1068
rect 8078 -1158 8112 -1124
rect 8146 -1158 8179 -1124
rect 8078 -1214 8179 -1158
rect 8078 -1248 8112 -1214
rect 8146 -1248 8179 -1214
rect 8078 -1304 8179 -1248
rect 9265 -348 9299 -314
rect 9333 -348 9366 -314
rect 9265 -404 9366 -348
rect 9265 -438 9299 -404
rect 9333 -438 9366 -404
rect 9265 -494 9366 -438
rect 9265 -528 9299 -494
rect 9333 -528 9366 -494
rect 9265 -584 9366 -528
rect 9265 -618 9299 -584
rect 9333 -618 9366 -584
rect 9265 -674 9366 -618
rect 9265 -708 9299 -674
rect 9333 -708 9366 -674
rect 9265 -764 9366 -708
rect 9265 -798 9299 -764
rect 9333 -798 9366 -764
rect 9265 -854 9366 -798
rect 9265 -888 9299 -854
rect 9333 -888 9366 -854
rect 9265 -944 9366 -888
rect 9265 -978 9299 -944
rect 9333 -978 9366 -944
rect 9265 -1034 9366 -978
rect 9265 -1068 9299 -1034
rect 9333 -1068 9366 -1034
rect 9265 -1124 9366 -1068
rect 9265 -1158 9299 -1124
rect 9333 -1158 9366 -1124
rect 9265 -1214 9366 -1158
rect 9265 -1248 9299 -1214
rect 9333 -1248 9366 -1214
rect 8078 -1338 8112 -1304
rect 8146 -1338 8179 -1304
rect 8078 -1353 8179 -1338
rect 9265 -1304 9366 -1248
rect 9265 -1338 9299 -1304
rect 9333 -1338 9366 -1304
rect 9265 -1353 9366 -1338
rect 8078 -1388 9366 -1353
rect 8078 -1422 8208 -1388
rect 8242 -1422 8298 -1388
rect 8332 -1422 8388 -1388
rect 8422 -1422 8478 -1388
rect 8512 -1422 8568 -1388
rect 8602 -1422 8658 -1388
rect 8692 -1422 8748 -1388
rect 8782 -1422 8838 -1388
rect 8872 -1422 8928 -1388
rect 8962 -1422 9018 -1388
rect 9052 -1422 9108 -1388
rect 9142 -1422 9198 -1388
rect 9232 -1422 9366 -1388
rect 8078 -1454 9366 -1422
<< nsubdiff >>
rect 189 3678 1151 3697
rect 189 3644 320 3678
rect 354 3644 410 3678
rect 444 3644 500 3678
rect 534 3644 590 3678
rect 624 3644 680 3678
rect 714 3644 770 3678
rect 804 3644 860 3678
rect 894 3644 950 3678
rect 984 3644 1040 3678
rect 1074 3644 1151 3678
rect 189 3625 1151 3644
rect 189 3621 261 3625
rect 189 3587 208 3621
rect 242 3587 261 3621
rect 189 3531 261 3587
rect 1079 3602 1151 3625
rect 1079 3568 1098 3602
rect 1132 3568 1151 3602
rect 189 3497 208 3531
rect 242 3497 261 3531
rect 189 3441 261 3497
rect 189 3407 208 3441
rect 242 3407 261 3441
rect 189 3351 261 3407
rect 189 3317 208 3351
rect 242 3317 261 3351
rect 189 3261 261 3317
rect 189 3227 208 3261
rect 242 3227 261 3261
rect 189 3171 261 3227
rect 189 3137 208 3171
rect 242 3137 261 3171
rect 189 3081 261 3137
rect 189 3047 208 3081
rect 242 3047 261 3081
rect 189 2991 261 3047
rect 189 2957 208 2991
rect 242 2957 261 2991
rect 189 2901 261 2957
rect 189 2867 208 2901
rect 242 2867 261 2901
rect 1079 3512 1151 3568
rect 1079 3478 1098 3512
rect 1132 3478 1151 3512
rect 1079 3422 1151 3478
rect 1079 3388 1098 3422
rect 1132 3388 1151 3422
rect 1079 3332 1151 3388
rect 1079 3298 1098 3332
rect 1132 3298 1151 3332
rect 1079 3242 1151 3298
rect 1079 3208 1098 3242
rect 1132 3208 1151 3242
rect 1079 3152 1151 3208
rect 1079 3118 1098 3152
rect 1132 3118 1151 3152
rect 1079 3062 1151 3118
rect 1079 3028 1098 3062
rect 1132 3028 1151 3062
rect 1079 2972 1151 3028
rect 1079 2938 1098 2972
rect 1132 2938 1151 2972
rect 1079 2882 1151 2938
rect 189 2807 261 2867
rect 1079 2848 1098 2882
rect 1132 2848 1151 2882
rect 1079 2807 1151 2848
rect 189 2788 1151 2807
rect 189 2754 286 2788
rect 320 2754 376 2788
rect 410 2754 466 2788
rect 500 2754 556 2788
rect 590 2754 646 2788
rect 680 2754 736 2788
rect 770 2754 826 2788
rect 860 2754 916 2788
rect 950 2754 1006 2788
rect 1040 2754 1151 2788
rect 189 2735 1151 2754
rect 1531 3678 2493 3697
rect 1531 3644 1662 3678
rect 1696 3644 1752 3678
rect 1786 3644 1842 3678
rect 1876 3644 1932 3678
rect 1966 3644 2022 3678
rect 2056 3644 2112 3678
rect 2146 3644 2202 3678
rect 2236 3644 2292 3678
rect 2326 3644 2382 3678
rect 2416 3644 2493 3678
rect 1531 3625 2493 3644
rect 1531 3621 1603 3625
rect 1531 3587 1550 3621
rect 1584 3587 1603 3621
rect 1531 3531 1603 3587
rect 2421 3602 2493 3625
rect 2421 3568 2440 3602
rect 2474 3568 2493 3602
rect 1531 3497 1550 3531
rect 1584 3497 1603 3531
rect 1531 3441 1603 3497
rect 1531 3407 1550 3441
rect 1584 3407 1603 3441
rect 1531 3351 1603 3407
rect 1531 3317 1550 3351
rect 1584 3317 1603 3351
rect 1531 3261 1603 3317
rect 1531 3227 1550 3261
rect 1584 3227 1603 3261
rect 1531 3171 1603 3227
rect 1531 3137 1550 3171
rect 1584 3137 1603 3171
rect 1531 3081 1603 3137
rect 1531 3047 1550 3081
rect 1584 3047 1603 3081
rect 1531 2991 1603 3047
rect 1531 2957 1550 2991
rect 1584 2957 1603 2991
rect 1531 2901 1603 2957
rect 1531 2867 1550 2901
rect 1584 2867 1603 2901
rect 2421 3512 2493 3568
rect 2421 3478 2440 3512
rect 2474 3478 2493 3512
rect 2421 3422 2493 3478
rect 2421 3388 2440 3422
rect 2474 3388 2493 3422
rect 2421 3332 2493 3388
rect 2421 3298 2440 3332
rect 2474 3298 2493 3332
rect 2421 3242 2493 3298
rect 2421 3208 2440 3242
rect 2474 3208 2493 3242
rect 2421 3152 2493 3208
rect 2421 3118 2440 3152
rect 2474 3118 2493 3152
rect 2421 3062 2493 3118
rect 2421 3028 2440 3062
rect 2474 3028 2493 3062
rect 2421 2972 2493 3028
rect 2421 2938 2440 2972
rect 2474 2938 2493 2972
rect 2421 2882 2493 2938
rect 1531 2807 1603 2867
rect 2421 2848 2440 2882
rect 2474 2848 2493 2882
rect 2421 2807 2493 2848
rect 1531 2788 2493 2807
rect 1531 2754 1628 2788
rect 1662 2754 1718 2788
rect 1752 2754 1808 2788
rect 1842 2754 1898 2788
rect 1932 2754 1988 2788
rect 2022 2754 2078 2788
rect 2112 2754 2168 2788
rect 2202 2754 2258 2788
rect 2292 2754 2348 2788
rect 2382 2754 2493 2788
rect 1531 2735 2493 2754
rect 2873 3678 3835 3697
rect 2873 3644 3004 3678
rect 3038 3644 3094 3678
rect 3128 3644 3184 3678
rect 3218 3644 3274 3678
rect 3308 3644 3364 3678
rect 3398 3644 3454 3678
rect 3488 3644 3544 3678
rect 3578 3644 3634 3678
rect 3668 3644 3724 3678
rect 3758 3644 3835 3678
rect 2873 3625 3835 3644
rect 2873 3621 2945 3625
rect 2873 3587 2892 3621
rect 2926 3587 2945 3621
rect 2873 3531 2945 3587
rect 3763 3602 3835 3625
rect 3763 3568 3782 3602
rect 3816 3568 3835 3602
rect 2873 3497 2892 3531
rect 2926 3497 2945 3531
rect 2873 3441 2945 3497
rect 2873 3407 2892 3441
rect 2926 3407 2945 3441
rect 2873 3351 2945 3407
rect 2873 3317 2892 3351
rect 2926 3317 2945 3351
rect 2873 3261 2945 3317
rect 2873 3227 2892 3261
rect 2926 3227 2945 3261
rect 2873 3171 2945 3227
rect 2873 3137 2892 3171
rect 2926 3137 2945 3171
rect 2873 3081 2945 3137
rect 2873 3047 2892 3081
rect 2926 3047 2945 3081
rect 2873 2991 2945 3047
rect 2873 2957 2892 2991
rect 2926 2957 2945 2991
rect 2873 2901 2945 2957
rect 2873 2867 2892 2901
rect 2926 2867 2945 2901
rect 3763 3512 3835 3568
rect 3763 3478 3782 3512
rect 3816 3478 3835 3512
rect 3763 3422 3835 3478
rect 3763 3388 3782 3422
rect 3816 3388 3835 3422
rect 3763 3332 3835 3388
rect 3763 3298 3782 3332
rect 3816 3298 3835 3332
rect 3763 3242 3835 3298
rect 3763 3208 3782 3242
rect 3816 3208 3835 3242
rect 3763 3152 3835 3208
rect 3763 3118 3782 3152
rect 3816 3118 3835 3152
rect 3763 3062 3835 3118
rect 3763 3028 3782 3062
rect 3816 3028 3835 3062
rect 3763 2972 3835 3028
rect 3763 2938 3782 2972
rect 3816 2938 3835 2972
rect 3763 2882 3835 2938
rect 2873 2807 2945 2867
rect 3763 2848 3782 2882
rect 3816 2848 3835 2882
rect 3763 2807 3835 2848
rect 2873 2788 3835 2807
rect 2873 2754 2970 2788
rect 3004 2754 3060 2788
rect 3094 2754 3150 2788
rect 3184 2754 3240 2788
rect 3274 2754 3330 2788
rect 3364 2754 3420 2788
rect 3454 2754 3510 2788
rect 3544 2754 3600 2788
rect 3634 2754 3690 2788
rect 3724 2754 3835 2788
rect 2873 2735 3835 2754
rect 4215 3678 5177 3697
rect 4215 3644 4346 3678
rect 4380 3644 4436 3678
rect 4470 3644 4526 3678
rect 4560 3644 4616 3678
rect 4650 3644 4706 3678
rect 4740 3644 4796 3678
rect 4830 3644 4886 3678
rect 4920 3644 4976 3678
rect 5010 3644 5066 3678
rect 5100 3644 5177 3678
rect 4215 3625 5177 3644
rect 4215 3621 4287 3625
rect 4215 3587 4234 3621
rect 4268 3587 4287 3621
rect 4215 3531 4287 3587
rect 5105 3602 5177 3625
rect 5105 3568 5124 3602
rect 5158 3568 5177 3602
rect 4215 3497 4234 3531
rect 4268 3497 4287 3531
rect 4215 3441 4287 3497
rect 4215 3407 4234 3441
rect 4268 3407 4287 3441
rect 4215 3351 4287 3407
rect 4215 3317 4234 3351
rect 4268 3317 4287 3351
rect 4215 3261 4287 3317
rect 4215 3227 4234 3261
rect 4268 3227 4287 3261
rect 4215 3171 4287 3227
rect 4215 3137 4234 3171
rect 4268 3137 4287 3171
rect 4215 3081 4287 3137
rect 4215 3047 4234 3081
rect 4268 3047 4287 3081
rect 4215 2991 4287 3047
rect 4215 2957 4234 2991
rect 4268 2957 4287 2991
rect 4215 2901 4287 2957
rect 4215 2867 4234 2901
rect 4268 2867 4287 2901
rect 5105 3512 5177 3568
rect 5105 3478 5124 3512
rect 5158 3478 5177 3512
rect 5105 3422 5177 3478
rect 5105 3388 5124 3422
rect 5158 3388 5177 3422
rect 5105 3332 5177 3388
rect 5105 3298 5124 3332
rect 5158 3298 5177 3332
rect 5105 3242 5177 3298
rect 5105 3208 5124 3242
rect 5158 3208 5177 3242
rect 5105 3152 5177 3208
rect 5105 3118 5124 3152
rect 5158 3118 5177 3152
rect 5105 3062 5177 3118
rect 5105 3028 5124 3062
rect 5158 3028 5177 3062
rect 5105 2972 5177 3028
rect 5105 2938 5124 2972
rect 5158 2938 5177 2972
rect 5105 2882 5177 2938
rect 4215 2807 4287 2867
rect 5105 2848 5124 2882
rect 5158 2848 5177 2882
rect 5105 2807 5177 2848
rect 4215 2788 5177 2807
rect 4215 2754 4312 2788
rect 4346 2754 4402 2788
rect 4436 2754 4492 2788
rect 4526 2754 4582 2788
rect 4616 2754 4672 2788
rect 4706 2754 4762 2788
rect 4796 2754 4852 2788
rect 4886 2754 4942 2788
rect 4976 2754 5032 2788
rect 5066 2754 5177 2788
rect 4215 2735 5177 2754
rect 5557 3678 6519 3697
rect 5557 3644 5688 3678
rect 5722 3644 5778 3678
rect 5812 3644 5868 3678
rect 5902 3644 5958 3678
rect 5992 3644 6048 3678
rect 6082 3644 6138 3678
rect 6172 3644 6228 3678
rect 6262 3644 6318 3678
rect 6352 3644 6408 3678
rect 6442 3644 6519 3678
rect 5557 3625 6519 3644
rect 5557 3621 5629 3625
rect 5557 3587 5576 3621
rect 5610 3587 5629 3621
rect 5557 3531 5629 3587
rect 6447 3602 6519 3625
rect 6447 3568 6466 3602
rect 6500 3568 6519 3602
rect 5557 3497 5576 3531
rect 5610 3497 5629 3531
rect 5557 3441 5629 3497
rect 5557 3407 5576 3441
rect 5610 3407 5629 3441
rect 5557 3351 5629 3407
rect 5557 3317 5576 3351
rect 5610 3317 5629 3351
rect 5557 3261 5629 3317
rect 5557 3227 5576 3261
rect 5610 3227 5629 3261
rect 5557 3171 5629 3227
rect 5557 3137 5576 3171
rect 5610 3137 5629 3171
rect 5557 3081 5629 3137
rect 5557 3047 5576 3081
rect 5610 3047 5629 3081
rect 5557 2991 5629 3047
rect 5557 2957 5576 2991
rect 5610 2957 5629 2991
rect 5557 2901 5629 2957
rect 5557 2867 5576 2901
rect 5610 2867 5629 2901
rect 6447 3512 6519 3568
rect 6447 3478 6466 3512
rect 6500 3478 6519 3512
rect 6447 3422 6519 3478
rect 6447 3388 6466 3422
rect 6500 3388 6519 3422
rect 6447 3332 6519 3388
rect 6447 3298 6466 3332
rect 6500 3298 6519 3332
rect 6447 3242 6519 3298
rect 6447 3208 6466 3242
rect 6500 3208 6519 3242
rect 6447 3152 6519 3208
rect 6447 3118 6466 3152
rect 6500 3118 6519 3152
rect 6447 3062 6519 3118
rect 6447 3028 6466 3062
rect 6500 3028 6519 3062
rect 6447 2972 6519 3028
rect 6447 2938 6466 2972
rect 6500 2938 6519 2972
rect 6447 2882 6519 2938
rect 5557 2807 5629 2867
rect 6447 2848 6466 2882
rect 6500 2848 6519 2882
rect 6447 2807 6519 2848
rect 5557 2788 6519 2807
rect 5557 2754 5654 2788
rect 5688 2754 5744 2788
rect 5778 2754 5834 2788
rect 5868 2754 5924 2788
rect 5958 2754 6014 2788
rect 6048 2754 6104 2788
rect 6138 2754 6194 2788
rect 6228 2754 6284 2788
rect 6318 2754 6374 2788
rect 6408 2754 6519 2788
rect 5557 2735 6519 2754
rect 6899 3678 7861 3697
rect 6899 3644 7030 3678
rect 7064 3644 7120 3678
rect 7154 3644 7210 3678
rect 7244 3644 7300 3678
rect 7334 3644 7390 3678
rect 7424 3644 7480 3678
rect 7514 3644 7570 3678
rect 7604 3644 7660 3678
rect 7694 3644 7750 3678
rect 7784 3644 7861 3678
rect 6899 3625 7861 3644
rect 6899 3621 6971 3625
rect 6899 3587 6918 3621
rect 6952 3587 6971 3621
rect 6899 3531 6971 3587
rect 7789 3602 7861 3625
rect 7789 3568 7808 3602
rect 7842 3568 7861 3602
rect 6899 3497 6918 3531
rect 6952 3497 6971 3531
rect 6899 3441 6971 3497
rect 6899 3407 6918 3441
rect 6952 3407 6971 3441
rect 6899 3351 6971 3407
rect 6899 3317 6918 3351
rect 6952 3317 6971 3351
rect 6899 3261 6971 3317
rect 6899 3227 6918 3261
rect 6952 3227 6971 3261
rect 6899 3171 6971 3227
rect 6899 3137 6918 3171
rect 6952 3137 6971 3171
rect 6899 3081 6971 3137
rect 6899 3047 6918 3081
rect 6952 3047 6971 3081
rect 6899 2991 6971 3047
rect 6899 2957 6918 2991
rect 6952 2957 6971 2991
rect 6899 2901 6971 2957
rect 6899 2867 6918 2901
rect 6952 2867 6971 2901
rect 7789 3512 7861 3568
rect 7789 3478 7808 3512
rect 7842 3478 7861 3512
rect 7789 3422 7861 3478
rect 7789 3388 7808 3422
rect 7842 3388 7861 3422
rect 7789 3332 7861 3388
rect 7789 3298 7808 3332
rect 7842 3298 7861 3332
rect 7789 3242 7861 3298
rect 7789 3208 7808 3242
rect 7842 3208 7861 3242
rect 7789 3152 7861 3208
rect 7789 3118 7808 3152
rect 7842 3118 7861 3152
rect 7789 3062 7861 3118
rect 7789 3028 7808 3062
rect 7842 3028 7861 3062
rect 7789 2972 7861 3028
rect 7789 2938 7808 2972
rect 7842 2938 7861 2972
rect 7789 2882 7861 2938
rect 6899 2807 6971 2867
rect 7789 2848 7808 2882
rect 7842 2848 7861 2882
rect 7789 2807 7861 2848
rect 6899 2788 7861 2807
rect 6899 2754 6996 2788
rect 7030 2754 7086 2788
rect 7120 2754 7176 2788
rect 7210 2754 7266 2788
rect 7300 2754 7356 2788
rect 7390 2754 7446 2788
rect 7480 2754 7536 2788
rect 7570 2754 7626 2788
rect 7660 2754 7716 2788
rect 7750 2754 7861 2788
rect 6899 2735 7861 2754
rect 8241 3678 9203 3697
rect 8241 3644 8372 3678
rect 8406 3644 8462 3678
rect 8496 3644 8552 3678
rect 8586 3644 8642 3678
rect 8676 3644 8732 3678
rect 8766 3644 8822 3678
rect 8856 3644 8912 3678
rect 8946 3644 9002 3678
rect 9036 3644 9092 3678
rect 9126 3644 9203 3678
rect 8241 3625 9203 3644
rect 8241 3621 8313 3625
rect 8241 3587 8260 3621
rect 8294 3587 8313 3621
rect 8241 3531 8313 3587
rect 9131 3602 9203 3625
rect 9131 3568 9150 3602
rect 9184 3568 9203 3602
rect 8241 3497 8260 3531
rect 8294 3497 8313 3531
rect 8241 3441 8313 3497
rect 8241 3407 8260 3441
rect 8294 3407 8313 3441
rect 8241 3351 8313 3407
rect 8241 3317 8260 3351
rect 8294 3317 8313 3351
rect 8241 3261 8313 3317
rect 8241 3227 8260 3261
rect 8294 3227 8313 3261
rect 8241 3171 8313 3227
rect 8241 3137 8260 3171
rect 8294 3137 8313 3171
rect 8241 3081 8313 3137
rect 8241 3047 8260 3081
rect 8294 3047 8313 3081
rect 8241 2991 8313 3047
rect 8241 2957 8260 2991
rect 8294 2957 8313 2991
rect 8241 2901 8313 2957
rect 8241 2867 8260 2901
rect 8294 2867 8313 2901
rect 9131 3512 9203 3568
rect 9131 3478 9150 3512
rect 9184 3478 9203 3512
rect 9131 3422 9203 3478
rect 9131 3388 9150 3422
rect 9184 3388 9203 3422
rect 9131 3332 9203 3388
rect 9131 3298 9150 3332
rect 9184 3298 9203 3332
rect 9131 3242 9203 3298
rect 9131 3208 9150 3242
rect 9184 3208 9203 3242
rect 9131 3152 9203 3208
rect 9131 3118 9150 3152
rect 9184 3118 9203 3152
rect 9131 3062 9203 3118
rect 9131 3028 9150 3062
rect 9184 3028 9203 3062
rect 9131 2972 9203 3028
rect 9131 2938 9150 2972
rect 9184 2938 9203 2972
rect 9131 2882 9203 2938
rect 8241 2807 8313 2867
rect 9131 2848 9150 2882
rect 9184 2848 9203 2882
rect 9131 2807 9203 2848
rect 8241 2788 9203 2807
rect 8241 2754 8338 2788
rect 8372 2754 8428 2788
rect 8462 2754 8518 2788
rect 8552 2754 8608 2788
rect 8642 2754 8698 2788
rect 8732 2754 8788 2788
rect 8822 2754 8878 2788
rect 8912 2754 8968 2788
rect 9002 2754 9058 2788
rect 9092 2754 9203 2788
rect 8241 2735 9203 2754
rect 189 2336 1151 2355
rect 189 2302 320 2336
rect 354 2302 410 2336
rect 444 2302 500 2336
rect 534 2302 590 2336
rect 624 2302 680 2336
rect 714 2302 770 2336
rect 804 2302 860 2336
rect 894 2302 950 2336
rect 984 2302 1040 2336
rect 1074 2302 1151 2336
rect 189 2283 1151 2302
rect 189 2279 261 2283
rect 189 2245 208 2279
rect 242 2245 261 2279
rect 189 2189 261 2245
rect 1079 2260 1151 2283
rect 1079 2226 1098 2260
rect 1132 2226 1151 2260
rect 189 2155 208 2189
rect 242 2155 261 2189
rect 189 2099 261 2155
rect 189 2065 208 2099
rect 242 2065 261 2099
rect 189 2009 261 2065
rect 189 1975 208 2009
rect 242 1975 261 2009
rect 189 1919 261 1975
rect 189 1885 208 1919
rect 242 1885 261 1919
rect 189 1829 261 1885
rect 189 1795 208 1829
rect 242 1795 261 1829
rect 189 1739 261 1795
rect 189 1705 208 1739
rect 242 1705 261 1739
rect 189 1649 261 1705
rect 189 1615 208 1649
rect 242 1615 261 1649
rect 189 1559 261 1615
rect 189 1525 208 1559
rect 242 1525 261 1559
rect 1079 2170 1151 2226
rect 1079 2136 1098 2170
rect 1132 2136 1151 2170
rect 1079 2080 1151 2136
rect 1079 2046 1098 2080
rect 1132 2046 1151 2080
rect 1079 1990 1151 2046
rect 1079 1956 1098 1990
rect 1132 1956 1151 1990
rect 1079 1900 1151 1956
rect 1079 1866 1098 1900
rect 1132 1866 1151 1900
rect 1079 1810 1151 1866
rect 1079 1776 1098 1810
rect 1132 1776 1151 1810
rect 1079 1720 1151 1776
rect 1079 1686 1098 1720
rect 1132 1686 1151 1720
rect 1079 1630 1151 1686
rect 1079 1596 1098 1630
rect 1132 1596 1151 1630
rect 1079 1540 1151 1596
rect 189 1465 261 1525
rect 1079 1506 1098 1540
rect 1132 1506 1151 1540
rect 1079 1465 1151 1506
rect 189 1446 1151 1465
rect 189 1412 286 1446
rect 320 1412 376 1446
rect 410 1412 466 1446
rect 500 1412 556 1446
rect 590 1412 646 1446
rect 680 1412 736 1446
rect 770 1412 826 1446
rect 860 1412 916 1446
rect 950 1412 1006 1446
rect 1040 1412 1151 1446
rect 189 1393 1151 1412
rect 1531 2336 2493 2355
rect 1531 2302 1662 2336
rect 1696 2302 1752 2336
rect 1786 2302 1842 2336
rect 1876 2302 1932 2336
rect 1966 2302 2022 2336
rect 2056 2302 2112 2336
rect 2146 2302 2202 2336
rect 2236 2302 2292 2336
rect 2326 2302 2382 2336
rect 2416 2302 2493 2336
rect 1531 2283 2493 2302
rect 1531 2279 1603 2283
rect 1531 2245 1550 2279
rect 1584 2245 1603 2279
rect 1531 2189 1603 2245
rect 2421 2260 2493 2283
rect 2421 2226 2440 2260
rect 2474 2226 2493 2260
rect 1531 2155 1550 2189
rect 1584 2155 1603 2189
rect 1531 2099 1603 2155
rect 1531 2065 1550 2099
rect 1584 2065 1603 2099
rect 1531 2009 1603 2065
rect 1531 1975 1550 2009
rect 1584 1975 1603 2009
rect 1531 1919 1603 1975
rect 1531 1885 1550 1919
rect 1584 1885 1603 1919
rect 1531 1829 1603 1885
rect 1531 1795 1550 1829
rect 1584 1795 1603 1829
rect 1531 1739 1603 1795
rect 1531 1705 1550 1739
rect 1584 1705 1603 1739
rect 1531 1649 1603 1705
rect 1531 1615 1550 1649
rect 1584 1615 1603 1649
rect 1531 1559 1603 1615
rect 1531 1525 1550 1559
rect 1584 1525 1603 1559
rect 2421 2170 2493 2226
rect 2421 2136 2440 2170
rect 2474 2136 2493 2170
rect 2421 2080 2493 2136
rect 2421 2046 2440 2080
rect 2474 2046 2493 2080
rect 2421 1990 2493 2046
rect 2421 1956 2440 1990
rect 2474 1956 2493 1990
rect 2421 1900 2493 1956
rect 2421 1866 2440 1900
rect 2474 1866 2493 1900
rect 2421 1810 2493 1866
rect 2421 1776 2440 1810
rect 2474 1776 2493 1810
rect 2421 1720 2493 1776
rect 2421 1686 2440 1720
rect 2474 1686 2493 1720
rect 2421 1630 2493 1686
rect 2421 1596 2440 1630
rect 2474 1596 2493 1630
rect 2421 1540 2493 1596
rect 1531 1465 1603 1525
rect 2421 1506 2440 1540
rect 2474 1506 2493 1540
rect 2421 1465 2493 1506
rect 1531 1446 2493 1465
rect 1531 1412 1628 1446
rect 1662 1412 1718 1446
rect 1752 1412 1808 1446
rect 1842 1412 1898 1446
rect 1932 1412 1988 1446
rect 2022 1412 2078 1446
rect 2112 1412 2168 1446
rect 2202 1412 2258 1446
rect 2292 1412 2348 1446
rect 2382 1412 2493 1446
rect 1531 1393 2493 1412
rect 2873 2336 3835 2355
rect 2873 2302 3004 2336
rect 3038 2302 3094 2336
rect 3128 2302 3184 2336
rect 3218 2302 3274 2336
rect 3308 2302 3364 2336
rect 3398 2302 3454 2336
rect 3488 2302 3544 2336
rect 3578 2302 3634 2336
rect 3668 2302 3724 2336
rect 3758 2302 3835 2336
rect 2873 2283 3835 2302
rect 2873 2279 2945 2283
rect 2873 2245 2892 2279
rect 2926 2245 2945 2279
rect 2873 2189 2945 2245
rect 3763 2260 3835 2283
rect 3763 2226 3782 2260
rect 3816 2226 3835 2260
rect 2873 2155 2892 2189
rect 2926 2155 2945 2189
rect 2873 2099 2945 2155
rect 2873 2065 2892 2099
rect 2926 2065 2945 2099
rect 2873 2009 2945 2065
rect 2873 1975 2892 2009
rect 2926 1975 2945 2009
rect 2873 1919 2945 1975
rect 2873 1885 2892 1919
rect 2926 1885 2945 1919
rect 2873 1829 2945 1885
rect 2873 1795 2892 1829
rect 2926 1795 2945 1829
rect 2873 1739 2945 1795
rect 2873 1705 2892 1739
rect 2926 1705 2945 1739
rect 2873 1649 2945 1705
rect 2873 1615 2892 1649
rect 2926 1615 2945 1649
rect 2873 1559 2945 1615
rect 2873 1525 2892 1559
rect 2926 1525 2945 1559
rect 3763 2170 3835 2226
rect 3763 2136 3782 2170
rect 3816 2136 3835 2170
rect 3763 2080 3835 2136
rect 3763 2046 3782 2080
rect 3816 2046 3835 2080
rect 3763 1990 3835 2046
rect 3763 1956 3782 1990
rect 3816 1956 3835 1990
rect 3763 1900 3835 1956
rect 3763 1866 3782 1900
rect 3816 1866 3835 1900
rect 3763 1810 3835 1866
rect 3763 1776 3782 1810
rect 3816 1776 3835 1810
rect 3763 1720 3835 1776
rect 3763 1686 3782 1720
rect 3816 1686 3835 1720
rect 3763 1630 3835 1686
rect 3763 1596 3782 1630
rect 3816 1596 3835 1630
rect 3763 1540 3835 1596
rect 2873 1465 2945 1525
rect 3763 1506 3782 1540
rect 3816 1506 3835 1540
rect 3763 1465 3835 1506
rect 2873 1446 3835 1465
rect 2873 1412 2970 1446
rect 3004 1412 3060 1446
rect 3094 1412 3150 1446
rect 3184 1412 3240 1446
rect 3274 1412 3330 1446
rect 3364 1412 3420 1446
rect 3454 1412 3510 1446
rect 3544 1412 3600 1446
rect 3634 1412 3690 1446
rect 3724 1412 3835 1446
rect 2873 1393 3835 1412
rect 4215 2336 5177 2355
rect 4215 2302 4346 2336
rect 4380 2302 4436 2336
rect 4470 2302 4526 2336
rect 4560 2302 4616 2336
rect 4650 2302 4706 2336
rect 4740 2302 4796 2336
rect 4830 2302 4886 2336
rect 4920 2302 4976 2336
rect 5010 2302 5066 2336
rect 5100 2302 5177 2336
rect 4215 2283 5177 2302
rect 4215 2279 4287 2283
rect 4215 2245 4234 2279
rect 4268 2245 4287 2279
rect 4215 2189 4287 2245
rect 5105 2260 5177 2283
rect 5105 2226 5124 2260
rect 5158 2226 5177 2260
rect 4215 2155 4234 2189
rect 4268 2155 4287 2189
rect 4215 2099 4287 2155
rect 4215 2065 4234 2099
rect 4268 2065 4287 2099
rect 4215 2009 4287 2065
rect 4215 1975 4234 2009
rect 4268 1975 4287 2009
rect 4215 1919 4287 1975
rect 4215 1885 4234 1919
rect 4268 1885 4287 1919
rect 4215 1829 4287 1885
rect 4215 1795 4234 1829
rect 4268 1795 4287 1829
rect 4215 1739 4287 1795
rect 4215 1705 4234 1739
rect 4268 1705 4287 1739
rect 4215 1649 4287 1705
rect 4215 1615 4234 1649
rect 4268 1615 4287 1649
rect 4215 1559 4287 1615
rect 4215 1525 4234 1559
rect 4268 1525 4287 1559
rect 5105 2170 5177 2226
rect 5105 2136 5124 2170
rect 5158 2136 5177 2170
rect 5105 2080 5177 2136
rect 5105 2046 5124 2080
rect 5158 2046 5177 2080
rect 5105 1990 5177 2046
rect 5105 1956 5124 1990
rect 5158 1956 5177 1990
rect 5105 1900 5177 1956
rect 5105 1866 5124 1900
rect 5158 1866 5177 1900
rect 5105 1810 5177 1866
rect 5105 1776 5124 1810
rect 5158 1776 5177 1810
rect 5105 1720 5177 1776
rect 5105 1686 5124 1720
rect 5158 1686 5177 1720
rect 5105 1630 5177 1686
rect 5105 1596 5124 1630
rect 5158 1596 5177 1630
rect 5105 1540 5177 1596
rect 4215 1465 4287 1525
rect 5105 1506 5124 1540
rect 5158 1506 5177 1540
rect 5105 1465 5177 1506
rect 4215 1446 5177 1465
rect 4215 1412 4312 1446
rect 4346 1412 4402 1446
rect 4436 1412 4492 1446
rect 4526 1412 4582 1446
rect 4616 1412 4672 1446
rect 4706 1412 4762 1446
rect 4796 1412 4852 1446
rect 4886 1412 4942 1446
rect 4976 1412 5032 1446
rect 5066 1412 5177 1446
rect 4215 1393 5177 1412
rect 5557 2336 6519 2355
rect 5557 2302 5688 2336
rect 5722 2302 5778 2336
rect 5812 2302 5868 2336
rect 5902 2302 5958 2336
rect 5992 2302 6048 2336
rect 6082 2302 6138 2336
rect 6172 2302 6228 2336
rect 6262 2302 6318 2336
rect 6352 2302 6408 2336
rect 6442 2302 6519 2336
rect 5557 2283 6519 2302
rect 5557 2279 5629 2283
rect 5557 2245 5576 2279
rect 5610 2245 5629 2279
rect 5557 2189 5629 2245
rect 6447 2260 6519 2283
rect 6447 2226 6466 2260
rect 6500 2226 6519 2260
rect 5557 2155 5576 2189
rect 5610 2155 5629 2189
rect 5557 2099 5629 2155
rect 5557 2065 5576 2099
rect 5610 2065 5629 2099
rect 5557 2009 5629 2065
rect 5557 1975 5576 2009
rect 5610 1975 5629 2009
rect 5557 1919 5629 1975
rect 5557 1885 5576 1919
rect 5610 1885 5629 1919
rect 5557 1829 5629 1885
rect 5557 1795 5576 1829
rect 5610 1795 5629 1829
rect 5557 1739 5629 1795
rect 5557 1705 5576 1739
rect 5610 1705 5629 1739
rect 5557 1649 5629 1705
rect 5557 1615 5576 1649
rect 5610 1615 5629 1649
rect 5557 1559 5629 1615
rect 5557 1525 5576 1559
rect 5610 1525 5629 1559
rect 6447 2170 6519 2226
rect 6447 2136 6466 2170
rect 6500 2136 6519 2170
rect 6447 2080 6519 2136
rect 6447 2046 6466 2080
rect 6500 2046 6519 2080
rect 6447 1990 6519 2046
rect 6447 1956 6466 1990
rect 6500 1956 6519 1990
rect 6447 1900 6519 1956
rect 6447 1866 6466 1900
rect 6500 1866 6519 1900
rect 6447 1810 6519 1866
rect 6447 1776 6466 1810
rect 6500 1776 6519 1810
rect 6447 1720 6519 1776
rect 6447 1686 6466 1720
rect 6500 1686 6519 1720
rect 6447 1630 6519 1686
rect 6447 1596 6466 1630
rect 6500 1596 6519 1630
rect 6447 1540 6519 1596
rect 5557 1465 5629 1525
rect 6447 1506 6466 1540
rect 6500 1506 6519 1540
rect 6447 1465 6519 1506
rect 5557 1446 6519 1465
rect 5557 1412 5654 1446
rect 5688 1412 5744 1446
rect 5778 1412 5834 1446
rect 5868 1412 5924 1446
rect 5958 1412 6014 1446
rect 6048 1412 6104 1446
rect 6138 1412 6194 1446
rect 6228 1412 6284 1446
rect 6318 1412 6374 1446
rect 6408 1412 6519 1446
rect 5557 1393 6519 1412
rect 6899 2336 7861 2355
rect 6899 2302 7030 2336
rect 7064 2302 7120 2336
rect 7154 2302 7210 2336
rect 7244 2302 7300 2336
rect 7334 2302 7390 2336
rect 7424 2302 7480 2336
rect 7514 2302 7570 2336
rect 7604 2302 7660 2336
rect 7694 2302 7750 2336
rect 7784 2302 7861 2336
rect 6899 2283 7861 2302
rect 6899 2279 6971 2283
rect 6899 2245 6918 2279
rect 6952 2245 6971 2279
rect 6899 2189 6971 2245
rect 7789 2260 7861 2283
rect 7789 2226 7808 2260
rect 7842 2226 7861 2260
rect 6899 2155 6918 2189
rect 6952 2155 6971 2189
rect 6899 2099 6971 2155
rect 6899 2065 6918 2099
rect 6952 2065 6971 2099
rect 6899 2009 6971 2065
rect 6899 1975 6918 2009
rect 6952 1975 6971 2009
rect 6899 1919 6971 1975
rect 6899 1885 6918 1919
rect 6952 1885 6971 1919
rect 6899 1829 6971 1885
rect 6899 1795 6918 1829
rect 6952 1795 6971 1829
rect 6899 1739 6971 1795
rect 6899 1705 6918 1739
rect 6952 1705 6971 1739
rect 6899 1649 6971 1705
rect 6899 1615 6918 1649
rect 6952 1615 6971 1649
rect 6899 1559 6971 1615
rect 6899 1525 6918 1559
rect 6952 1525 6971 1559
rect 7789 2170 7861 2226
rect 7789 2136 7808 2170
rect 7842 2136 7861 2170
rect 7789 2080 7861 2136
rect 7789 2046 7808 2080
rect 7842 2046 7861 2080
rect 7789 1990 7861 2046
rect 7789 1956 7808 1990
rect 7842 1956 7861 1990
rect 7789 1900 7861 1956
rect 7789 1866 7808 1900
rect 7842 1866 7861 1900
rect 7789 1810 7861 1866
rect 7789 1776 7808 1810
rect 7842 1776 7861 1810
rect 7789 1720 7861 1776
rect 7789 1686 7808 1720
rect 7842 1686 7861 1720
rect 7789 1630 7861 1686
rect 7789 1596 7808 1630
rect 7842 1596 7861 1630
rect 7789 1540 7861 1596
rect 6899 1465 6971 1525
rect 7789 1506 7808 1540
rect 7842 1506 7861 1540
rect 7789 1465 7861 1506
rect 6899 1446 7861 1465
rect 6899 1412 6996 1446
rect 7030 1412 7086 1446
rect 7120 1412 7176 1446
rect 7210 1412 7266 1446
rect 7300 1412 7356 1446
rect 7390 1412 7446 1446
rect 7480 1412 7536 1446
rect 7570 1412 7626 1446
rect 7660 1412 7716 1446
rect 7750 1412 7861 1446
rect 6899 1393 7861 1412
rect 8241 2336 9203 2355
rect 8241 2302 8372 2336
rect 8406 2302 8462 2336
rect 8496 2302 8552 2336
rect 8586 2302 8642 2336
rect 8676 2302 8732 2336
rect 8766 2302 8822 2336
rect 8856 2302 8912 2336
rect 8946 2302 9002 2336
rect 9036 2302 9092 2336
rect 9126 2302 9203 2336
rect 8241 2283 9203 2302
rect 8241 2279 8313 2283
rect 8241 2245 8260 2279
rect 8294 2245 8313 2279
rect 8241 2189 8313 2245
rect 9131 2260 9203 2283
rect 9131 2226 9150 2260
rect 9184 2226 9203 2260
rect 8241 2155 8260 2189
rect 8294 2155 8313 2189
rect 8241 2099 8313 2155
rect 8241 2065 8260 2099
rect 8294 2065 8313 2099
rect 8241 2009 8313 2065
rect 8241 1975 8260 2009
rect 8294 1975 8313 2009
rect 8241 1919 8313 1975
rect 8241 1885 8260 1919
rect 8294 1885 8313 1919
rect 8241 1829 8313 1885
rect 8241 1795 8260 1829
rect 8294 1795 8313 1829
rect 8241 1739 8313 1795
rect 8241 1705 8260 1739
rect 8294 1705 8313 1739
rect 8241 1649 8313 1705
rect 8241 1615 8260 1649
rect 8294 1615 8313 1649
rect 8241 1559 8313 1615
rect 8241 1525 8260 1559
rect 8294 1525 8313 1559
rect 9131 2170 9203 2226
rect 9131 2136 9150 2170
rect 9184 2136 9203 2170
rect 9131 2080 9203 2136
rect 9131 2046 9150 2080
rect 9184 2046 9203 2080
rect 9131 1990 9203 2046
rect 9131 1956 9150 1990
rect 9184 1956 9203 1990
rect 9131 1900 9203 1956
rect 9131 1866 9150 1900
rect 9184 1866 9203 1900
rect 9131 1810 9203 1866
rect 9131 1776 9150 1810
rect 9184 1776 9203 1810
rect 9131 1720 9203 1776
rect 9131 1686 9150 1720
rect 9184 1686 9203 1720
rect 9131 1630 9203 1686
rect 9131 1596 9150 1630
rect 9184 1596 9203 1630
rect 9131 1540 9203 1596
rect 8241 1465 8313 1525
rect 9131 1506 9150 1540
rect 9184 1506 9203 1540
rect 9131 1465 9203 1506
rect 8241 1446 9203 1465
rect 8241 1412 8338 1446
rect 8372 1412 8428 1446
rect 8462 1412 8518 1446
rect 8552 1412 8608 1446
rect 8642 1412 8698 1446
rect 8732 1412 8788 1446
rect 8822 1412 8878 1446
rect 8912 1412 8968 1446
rect 9002 1412 9058 1446
rect 9092 1412 9203 1446
rect 8241 1393 9203 1412
rect 1686 941 2493 1013
rect 1531 123 1603 874
rect 2421 123 2493 941
rect 1531 51 2493 123
rect 2873 941 3835 1013
rect 2873 123 2945 941
rect 3763 123 3835 941
rect 2873 51 3835 123
rect 4215 941 5177 1013
rect 4215 123 4287 941
rect 5105 123 5177 941
rect 4215 51 5177 123
rect 5557 941 6519 1013
rect 5557 123 5629 941
rect 6447 123 6519 941
rect 5557 51 6519 123
rect 6899 994 7861 1013
rect 6899 960 7030 994
rect 7064 960 7120 994
rect 7154 960 7210 994
rect 7244 960 7300 994
rect 7334 960 7390 994
rect 7424 960 7480 994
rect 7514 960 7570 994
rect 7604 960 7660 994
rect 7694 960 7750 994
rect 7784 960 7861 994
rect 6899 941 7861 960
rect 6899 937 6971 941
rect 6899 903 6918 937
rect 6952 903 6971 937
rect 6899 847 6971 903
rect 7789 918 7861 941
rect 7789 884 7808 918
rect 7842 884 7861 918
rect 6899 813 6918 847
rect 6952 813 6971 847
rect 6899 757 6971 813
rect 6899 723 6918 757
rect 6952 723 6971 757
rect 6899 667 6971 723
rect 6899 633 6918 667
rect 6952 633 6971 667
rect 6899 577 6971 633
rect 6899 543 6918 577
rect 6952 543 6971 577
rect 6899 487 6971 543
rect 6899 453 6918 487
rect 6952 453 6971 487
rect 6899 397 6971 453
rect 6899 363 6918 397
rect 6952 363 6971 397
rect 6899 307 6971 363
rect 6899 273 6918 307
rect 6952 273 6971 307
rect 6899 217 6971 273
rect 6899 183 6918 217
rect 6952 183 6971 217
rect 7789 828 7861 884
rect 7789 794 7808 828
rect 7842 794 7861 828
rect 7789 738 7861 794
rect 7789 704 7808 738
rect 7842 704 7861 738
rect 7789 648 7861 704
rect 7789 614 7808 648
rect 7842 614 7861 648
rect 7789 558 7861 614
rect 7789 524 7808 558
rect 7842 524 7861 558
rect 7789 468 7861 524
rect 7789 434 7808 468
rect 7842 434 7861 468
rect 7789 378 7861 434
rect 7789 344 7808 378
rect 7842 344 7861 378
rect 7789 288 7861 344
rect 7789 254 7808 288
rect 7842 254 7861 288
rect 7789 198 7861 254
rect 6899 123 6971 183
rect 7789 164 7808 198
rect 7842 164 7861 198
rect 7789 123 7861 164
rect 6899 104 7861 123
rect 6899 70 6996 104
rect 7030 70 7086 104
rect 7120 70 7176 104
rect 7210 70 7266 104
rect 7300 70 7356 104
rect 7390 70 7446 104
rect 7480 70 7536 104
rect 7570 70 7626 104
rect 7660 70 7716 104
rect 7750 70 7861 104
rect 6899 51 7861 70
rect 8241 994 9203 1013
rect 8241 960 8372 994
rect 8406 960 8462 994
rect 8496 960 8552 994
rect 8586 960 8642 994
rect 8676 960 8732 994
rect 8766 960 8822 994
rect 8856 960 8912 994
rect 8946 960 9002 994
rect 9036 960 9092 994
rect 9126 960 9203 994
rect 8241 941 9203 960
rect 8241 937 8313 941
rect 8241 903 8260 937
rect 8294 903 8313 937
rect 8241 847 8313 903
rect 9131 918 9203 941
rect 9131 884 9150 918
rect 9184 884 9203 918
rect 8241 813 8260 847
rect 8294 813 8313 847
rect 8241 757 8313 813
rect 8241 723 8260 757
rect 8294 723 8313 757
rect 8241 667 8313 723
rect 8241 633 8260 667
rect 8294 633 8313 667
rect 8241 577 8313 633
rect 8241 543 8260 577
rect 8294 543 8313 577
rect 8241 487 8313 543
rect 8241 453 8260 487
rect 8294 453 8313 487
rect 8241 397 8313 453
rect 8241 363 8260 397
rect 8294 363 8313 397
rect 8241 307 8313 363
rect 8241 273 8260 307
rect 8294 273 8313 307
rect 8241 217 8313 273
rect 8241 183 8260 217
rect 8294 183 8313 217
rect 9131 828 9203 884
rect 9131 794 9150 828
rect 9184 794 9203 828
rect 9131 738 9203 794
rect 9131 704 9150 738
rect 9184 704 9203 738
rect 9131 648 9203 704
rect 9131 614 9150 648
rect 9184 614 9203 648
rect 9131 558 9203 614
rect 9131 524 9150 558
rect 9184 524 9203 558
rect 9131 468 9203 524
rect 9131 434 9150 468
rect 9184 434 9203 468
rect 9131 378 9203 434
rect 9131 344 9150 378
rect 9184 344 9203 378
rect 9131 288 9203 344
rect 9131 254 9150 288
rect 9184 254 9203 288
rect 9131 198 9203 254
rect 8241 123 8313 183
rect 9131 164 9150 198
rect 9184 164 9203 198
rect 9131 123 9203 164
rect 8241 104 9203 123
rect 8241 70 8338 104
rect 8372 70 8428 104
rect 8462 70 8518 104
rect 8552 70 8608 104
rect 8642 70 8698 104
rect 8732 70 8788 104
rect 8822 70 8878 104
rect 8912 70 8968 104
rect 9002 70 9058 104
rect 9092 70 9203 104
rect 8241 51 9203 70
rect 189 -401 1151 -329
rect 189 -1219 261 -401
rect 1079 -1219 1151 -401
rect 189 -1291 1151 -1219
rect 1531 -401 2493 -329
rect 1531 -1219 1603 -401
rect 2421 -1219 2493 -401
rect 1531 -1291 2493 -1219
rect 2873 -401 3835 -329
rect 2873 -1219 2945 -401
rect 3763 -1219 3835 -401
rect 2873 -1291 3835 -1219
rect 4215 -401 5177 -329
rect 4215 -1219 4287 -401
rect 5105 -1219 5177 -401
rect 4215 -1291 5177 -1219
rect 5557 -401 6519 -329
rect 5557 -1219 5629 -401
rect 6447 -1219 6519 -401
rect 5557 -1291 6519 -1219
rect 6899 -348 7861 -329
rect 6899 -382 7030 -348
rect 7064 -382 7120 -348
rect 7154 -382 7210 -348
rect 7244 -382 7300 -348
rect 7334 -382 7390 -348
rect 7424 -382 7480 -348
rect 7514 -382 7570 -348
rect 7604 -382 7660 -348
rect 7694 -382 7750 -348
rect 7784 -382 7861 -348
rect 6899 -401 7861 -382
rect 6899 -405 6971 -401
rect 6899 -439 6918 -405
rect 6952 -439 6971 -405
rect 6899 -495 6971 -439
rect 7789 -424 7861 -401
rect 7789 -458 7808 -424
rect 7842 -458 7861 -424
rect 6899 -529 6918 -495
rect 6952 -529 6971 -495
rect 6899 -585 6971 -529
rect 6899 -619 6918 -585
rect 6952 -619 6971 -585
rect 6899 -675 6971 -619
rect 6899 -709 6918 -675
rect 6952 -709 6971 -675
rect 6899 -765 6971 -709
rect 6899 -799 6918 -765
rect 6952 -799 6971 -765
rect 6899 -855 6971 -799
rect 6899 -889 6918 -855
rect 6952 -889 6971 -855
rect 6899 -945 6971 -889
rect 6899 -979 6918 -945
rect 6952 -979 6971 -945
rect 6899 -1035 6971 -979
rect 6899 -1069 6918 -1035
rect 6952 -1069 6971 -1035
rect 6899 -1125 6971 -1069
rect 6899 -1159 6918 -1125
rect 6952 -1159 6971 -1125
rect 7789 -514 7861 -458
rect 7789 -548 7808 -514
rect 7842 -548 7861 -514
rect 7789 -604 7861 -548
rect 7789 -638 7808 -604
rect 7842 -638 7861 -604
rect 7789 -694 7861 -638
rect 7789 -728 7808 -694
rect 7842 -728 7861 -694
rect 7789 -784 7861 -728
rect 7789 -818 7808 -784
rect 7842 -818 7861 -784
rect 7789 -874 7861 -818
rect 7789 -908 7808 -874
rect 7842 -908 7861 -874
rect 7789 -964 7861 -908
rect 7789 -998 7808 -964
rect 7842 -998 7861 -964
rect 7789 -1054 7861 -998
rect 7789 -1088 7808 -1054
rect 7842 -1088 7861 -1054
rect 7789 -1144 7861 -1088
rect 6899 -1219 6971 -1159
rect 7789 -1178 7808 -1144
rect 7842 -1178 7861 -1144
rect 7789 -1219 7861 -1178
rect 6899 -1238 7861 -1219
rect 6899 -1272 6996 -1238
rect 7030 -1272 7086 -1238
rect 7120 -1272 7176 -1238
rect 7210 -1272 7266 -1238
rect 7300 -1272 7356 -1238
rect 7390 -1272 7446 -1238
rect 7480 -1272 7536 -1238
rect 7570 -1272 7626 -1238
rect 7660 -1272 7716 -1238
rect 7750 -1272 7861 -1238
rect 6899 -1291 7861 -1272
rect 8241 -348 9203 -329
rect 8241 -382 8372 -348
rect 8406 -382 8462 -348
rect 8496 -382 8552 -348
rect 8586 -382 8642 -348
rect 8676 -382 8732 -348
rect 8766 -382 8822 -348
rect 8856 -382 8912 -348
rect 8946 -382 9002 -348
rect 9036 -382 9092 -348
rect 9126 -382 9203 -348
rect 8241 -401 9203 -382
rect 8241 -405 8313 -401
rect 8241 -439 8260 -405
rect 8294 -439 8313 -405
rect 8241 -495 8313 -439
rect 9131 -424 9203 -401
rect 9131 -458 9150 -424
rect 9184 -458 9203 -424
rect 8241 -529 8260 -495
rect 8294 -529 8313 -495
rect 8241 -585 8313 -529
rect 8241 -619 8260 -585
rect 8294 -619 8313 -585
rect 8241 -675 8313 -619
rect 8241 -709 8260 -675
rect 8294 -709 8313 -675
rect 8241 -765 8313 -709
rect 8241 -799 8260 -765
rect 8294 -799 8313 -765
rect 8241 -855 8313 -799
rect 8241 -889 8260 -855
rect 8294 -889 8313 -855
rect 8241 -945 8313 -889
rect 8241 -979 8260 -945
rect 8294 -979 8313 -945
rect 8241 -1035 8313 -979
rect 8241 -1069 8260 -1035
rect 8294 -1069 8313 -1035
rect 8241 -1125 8313 -1069
rect 8241 -1159 8260 -1125
rect 8294 -1159 8313 -1125
rect 9131 -514 9203 -458
rect 9131 -548 9150 -514
rect 9184 -548 9203 -514
rect 9131 -604 9203 -548
rect 9131 -638 9150 -604
rect 9184 -638 9203 -604
rect 9131 -694 9203 -638
rect 9131 -728 9150 -694
rect 9184 -728 9203 -694
rect 9131 -784 9203 -728
rect 9131 -818 9150 -784
rect 9184 -818 9203 -784
rect 9131 -874 9203 -818
rect 9131 -908 9150 -874
rect 9184 -908 9203 -874
rect 9131 -964 9203 -908
rect 9131 -998 9150 -964
rect 9184 -998 9203 -964
rect 9131 -1054 9203 -998
rect 9131 -1088 9150 -1054
rect 9184 -1088 9203 -1054
rect 9131 -1144 9203 -1088
rect 8241 -1219 8313 -1159
rect 9131 -1178 9150 -1144
rect 9184 -1178 9203 -1144
rect 9131 -1219 9203 -1178
rect 8241 -1238 9203 -1219
rect 8241 -1272 8338 -1238
rect 8372 -1272 8428 -1238
rect 8462 -1272 8518 -1238
rect 8552 -1272 8608 -1238
rect 8642 -1272 8698 -1238
rect 8732 -1272 8788 -1238
rect 8822 -1272 8878 -1238
rect 8912 -1272 8968 -1238
rect 9002 -1272 9058 -1238
rect 9092 -1272 9203 -1238
rect 8241 -1291 9203 -1272
<< psubdiffcont >>
rect 60 3768 94 3802
rect 156 3791 190 3825
rect 246 3791 280 3825
rect 336 3791 370 3825
rect 426 3791 460 3825
rect 516 3791 550 3825
rect 606 3791 640 3825
rect 696 3791 730 3825
rect 786 3791 820 3825
rect 876 3791 910 3825
rect 966 3791 1000 3825
rect 1056 3791 1090 3825
rect 1146 3791 1180 3825
rect 1247 3768 1281 3802
rect 60 3678 94 3712
rect 60 3588 94 3622
rect 60 3498 94 3532
rect 60 3408 94 3442
rect 60 3318 94 3352
rect 60 3228 94 3262
rect 60 3138 94 3172
rect 60 3048 94 3082
rect 60 2958 94 2992
rect 60 2868 94 2902
rect 60 2778 94 2812
rect 1247 3678 1281 3712
rect 1247 3588 1281 3622
rect 1247 3498 1281 3532
rect 1247 3408 1281 3442
rect 1247 3318 1281 3352
rect 1247 3228 1281 3262
rect 1247 3138 1281 3172
rect 1247 3048 1281 3082
rect 1247 2958 1281 2992
rect 1247 2868 1281 2902
rect 1247 2778 1281 2812
rect 60 2688 94 2722
rect 1247 2688 1281 2722
rect 156 2604 190 2638
rect 246 2604 280 2638
rect 336 2604 370 2638
rect 426 2604 460 2638
rect 516 2604 550 2638
rect 606 2604 640 2638
rect 696 2604 730 2638
rect 786 2604 820 2638
rect 876 2604 910 2638
rect 966 2604 1000 2638
rect 1056 2604 1090 2638
rect 1146 2604 1180 2638
rect 1402 3768 1436 3802
rect 1498 3791 1532 3825
rect 1588 3791 1622 3825
rect 1678 3791 1712 3825
rect 1768 3791 1802 3825
rect 1858 3791 1892 3825
rect 1948 3791 1982 3825
rect 2038 3791 2072 3825
rect 2128 3791 2162 3825
rect 2218 3791 2252 3825
rect 2308 3791 2342 3825
rect 2398 3791 2432 3825
rect 2488 3791 2522 3825
rect 2589 3768 2623 3802
rect 1402 3678 1436 3712
rect 1402 3588 1436 3622
rect 1402 3498 1436 3532
rect 1402 3408 1436 3442
rect 1402 3318 1436 3352
rect 1402 3228 1436 3262
rect 1402 3138 1436 3172
rect 1402 3048 1436 3082
rect 1402 2958 1436 2992
rect 1402 2868 1436 2902
rect 1402 2778 1436 2812
rect 2589 3678 2623 3712
rect 2589 3588 2623 3622
rect 2589 3498 2623 3532
rect 2589 3408 2623 3442
rect 2589 3318 2623 3352
rect 2589 3228 2623 3262
rect 2589 3138 2623 3172
rect 2589 3048 2623 3082
rect 2589 2958 2623 2992
rect 2589 2868 2623 2902
rect 2589 2778 2623 2812
rect 1402 2688 1436 2722
rect 2589 2688 2623 2722
rect 1498 2604 1532 2638
rect 1588 2604 1622 2638
rect 1678 2604 1712 2638
rect 1768 2604 1802 2638
rect 1858 2604 1892 2638
rect 1948 2604 1982 2638
rect 2038 2604 2072 2638
rect 2128 2604 2162 2638
rect 2218 2604 2252 2638
rect 2308 2604 2342 2638
rect 2398 2604 2432 2638
rect 2488 2604 2522 2638
rect 2744 3768 2778 3802
rect 2840 3791 2874 3825
rect 2930 3791 2964 3825
rect 3020 3791 3054 3825
rect 3110 3791 3144 3825
rect 3200 3791 3234 3825
rect 3290 3791 3324 3825
rect 3380 3791 3414 3825
rect 3470 3791 3504 3825
rect 3560 3791 3594 3825
rect 3650 3791 3684 3825
rect 3740 3791 3774 3825
rect 3830 3791 3864 3825
rect 3931 3768 3965 3802
rect 2744 3678 2778 3712
rect 2744 3588 2778 3622
rect 2744 3498 2778 3532
rect 2744 3408 2778 3442
rect 2744 3318 2778 3352
rect 2744 3228 2778 3262
rect 2744 3138 2778 3172
rect 2744 3048 2778 3082
rect 2744 2958 2778 2992
rect 2744 2868 2778 2902
rect 2744 2778 2778 2812
rect 3931 3678 3965 3712
rect 3931 3588 3965 3622
rect 3931 3498 3965 3532
rect 3931 3408 3965 3442
rect 3931 3318 3965 3352
rect 3931 3228 3965 3262
rect 3931 3138 3965 3172
rect 3931 3048 3965 3082
rect 3931 2958 3965 2992
rect 3931 2868 3965 2902
rect 3931 2778 3965 2812
rect 2744 2688 2778 2722
rect 3931 2688 3965 2722
rect 2840 2604 2874 2638
rect 2930 2604 2964 2638
rect 3020 2604 3054 2638
rect 3110 2604 3144 2638
rect 3200 2604 3234 2638
rect 3290 2604 3324 2638
rect 3380 2604 3414 2638
rect 3470 2604 3504 2638
rect 3560 2604 3594 2638
rect 3650 2604 3684 2638
rect 3740 2604 3774 2638
rect 3830 2604 3864 2638
rect 4086 3768 4120 3802
rect 4182 3791 4216 3825
rect 4272 3791 4306 3825
rect 4362 3791 4396 3825
rect 4452 3791 4486 3825
rect 4542 3791 4576 3825
rect 4632 3791 4666 3825
rect 4722 3791 4756 3825
rect 4812 3791 4846 3825
rect 4902 3791 4936 3825
rect 4992 3791 5026 3825
rect 5082 3791 5116 3825
rect 5172 3791 5206 3825
rect 5273 3768 5307 3802
rect 4086 3678 4120 3712
rect 4086 3588 4120 3622
rect 4086 3498 4120 3532
rect 4086 3408 4120 3442
rect 4086 3318 4120 3352
rect 4086 3228 4120 3262
rect 4086 3138 4120 3172
rect 4086 3048 4120 3082
rect 4086 2958 4120 2992
rect 4086 2868 4120 2902
rect 4086 2778 4120 2812
rect 5273 3678 5307 3712
rect 5273 3588 5307 3622
rect 5273 3498 5307 3532
rect 5273 3408 5307 3442
rect 5273 3318 5307 3352
rect 5273 3228 5307 3262
rect 5273 3138 5307 3172
rect 5273 3048 5307 3082
rect 5273 2958 5307 2992
rect 5273 2868 5307 2902
rect 5273 2778 5307 2812
rect 4086 2688 4120 2722
rect 5273 2688 5307 2722
rect 4182 2604 4216 2638
rect 4272 2604 4306 2638
rect 4362 2604 4396 2638
rect 4452 2604 4486 2638
rect 4542 2604 4576 2638
rect 4632 2604 4666 2638
rect 4722 2604 4756 2638
rect 4812 2604 4846 2638
rect 4902 2604 4936 2638
rect 4992 2604 5026 2638
rect 5082 2604 5116 2638
rect 5172 2604 5206 2638
rect 5428 3768 5462 3802
rect 5524 3791 5558 3825
rect 5614 3791 5648 3825
rect 5704 3791 5738 3825
rect 5794 3791 5828 3825
rect 5884 3791 5918 3825
rect 5974 3791 6008 3825
rect 6064 3791 6098 3825
rect 6154 3791 6188 3825
rect 6244 3791 6278 3825
rect 6334 3791 6368 3825
rect 6424 3791 6458 3825
rect 6514 3791 6548 3825
rect 6615 3768 6649 3802
rect 5428 3678 5462 3712
rect 5428 3588 5462 3622
rect 5428 3498 5462 3532
rect 5428 3408 5462 3442
rect 5428 3318 5462 3352
rect 5428 3228 5462 3262
rect 5428 3138 5462 3172
rect 5428 3048 5462 3082
rect 5428 2958 5462 2992
rect 5428 2868 5462 2902
rect 5428 2778 5462 2812
rect 6615 3678 6649 3712
rect 6615 3588 6649 3622
rect 6615 3498 6649 3532
rect 6615 3408 6649 3442
rect 6615 3318 6649 3352
rect 6615 3228 6649 3262
rect 6615 3138 6649 3172
rect 6615 3048 6649 3082
rect 6615 2958 6649 2992
rect 6615 2868 6649 2902
rect 6615 2778 6649 2812
rect 5428 2688 5462 2722
rect 6615 2688 6649 2722
rect 5524 2604 5558 2638
rect 5614 2604 5648 2638
rect 5704 2604 5738 2638
rect 5794 2604 5828 2638
rect 5884 2604 5918 2638
rect 5974 2604 6008 2638
rect 6064 2604 6098 2638
rect 6154 2604 6188 2638
rect 6244 2604 6278 2638
rect 6334 2604 6368 2638
rect 6424 2604 6458 2638
rect 6514 2604 6548 2638
rect 6770 3768 6804 3802
rect 6866 3791 6900 3825
rect 6956 3791 6990 3825
rect 7046 3791 7080 3825
rect 7136 3791 7170 3825
rect 7226 3791 7260 3825
rect 7316 3791 7350 3825
rect 7406 3791 7440 3825
rect 7496 3791 7530 3825
rect 7586 3791 7620 3825
rect 7676 3791 7710 3825
rect 7766 3791 7800 3825
rect 7856 3791 7890 3825
rect 7957 3768 7991 3802
rect 6770 3678 6804 3712
rect 6770 3588 6804 3622
rect 6770 3498 6804 3532
rect 6770 3408 6804 3442
rect 6770 3318 6804 3352
rect 6770 3228 6804 3262
rect 6770 3138 6804 3172
rect 6770 3048 6804 3082
rect 6770 2958 6804 2992
rect 6770 2868 6804 2902
rect 6770 2778 6804 2812
rect 7957 3678 7991 3712
rect 7957 3588 7991 3622
rect 7957 3498 7991 3532
rect 7957 3408 7991 3442
rect 7957 3318 7991 3352
rect 7957 3228 7991 3262
rect 7957 3138 7991 3172
rect 7957 3048 7991 3082
rect 7957 2958 7991 2992
rect 7957 2868 7991 2902
rect 7957 2778 7991 2812
rect 6770 2688 6804 2722
rect 7957 2688 7991 2722
rect 6866 2604 6900 2638
rect 6956 2604 6990 2638
rect 7046 2604 7080 2638
rect 7136 2604 7170 2638
rect 7226 2604 7260 2638
rect 7316 2604 7350 2638
rect 7406 2604 7440 2638
rect 7496 2604 7530 2638
rect 7586 2604 7620 2638
rect 7676 2604 7710 2638
rect 7766 2604 7800 2638
rect 7856 2604 7890 2638
rect 8112 3768 8146 3802
rect 8208 3791 8242 3825
rect 8298 3791 8332 3825
rect 8388 3791 8422 3825
rect 8478 3791 8512 3825
rect 8568 3791 8602 3825
rect 8658 3791 8692 3825
rect 8748 3791 8782 3825
rect 8838 3791 8872 3825
rect 8928 3791 8962 3825
rect 9018 3791 9052 3825
rect 9108 3791 9142 3825
rect 9198 3791 9232 3825
rect 9299 3768 9333 3802
rect 8112 3678 8146 3712
rect 8112 3588 8146 3622
rect 8112 3498 8146 3532
rect 8112 3408 8146 3442
rect 8112 3318 8146 3352
rect 8112 3228 8146 3262
rect 8112 3138 8146 3172
rect 8112 3048 8146 3082
rect 8112 2958 8146 2992
rect 8112 2868 8146 2902
rect 8112 2778 8146 2812
rect 9299 3678 9333 3712
rect 9299 3588 9333 3622
rect 9299 3498 9333 3532
rect 9299 3408 9333 3442
rect 9299 3318 9333 3352
rect 9299 3228 9333 3262
rect 9299 3138 9333 3172
rect 9299 3048 9333 3082
rect 9299 2958 9333 2992
rect 9299 2868 9333 2902
rect 9299 2778 9333 2812
rect 8112 2688 8146 2722
rect 9299 2688 9333 2722
rect 8208 2604 8242 2638
rect 8298 2604 8332 2638
rect 8388 2604 8422 2638
rect 8478 2604 8512 2638
rect 8568 2604 8602 2638
rect 8658 2604 8692 2638
rect 8748 2604 8782 2638
rect 8838 2604 8872 2638
rect 8928 2604 8962 2638
rect 9018 2604 9052 2638
rect 9108 2604 9142 2638
rect 9198 2604 9232 2638
rect 60 2426 94 2460
rect 156 2449 190 2483
rect 246 2449 280 2483
rect 336 2449 370 2483
rect 426 2449 460 2483
rect 516 2449 550 2483
rect 606 2449 640 2483
rect 696 2449 730 2483
rect 786 2449 820 2483
rect 876 2449 910 2483
rect 966 2449 1000 2483
rect 1056 2449 1090 2483
rect 1146 2449 1180 2483
rect 1247 2426 1281 2460
rect 60 2336 94 2370
rect 60 2246 94 2280
rect 60 2156 94 2190
rect 60 2066 94 2100
rect 60 1976 94 2010
rect 60 1886 94 1920
rect 60 1796 94 1830
rect 60 1706 94 1740
rect 60 1616 94 1650
rect 60 1526 94 1560
rect 60 1436 94 1470
rect 1247 2336 1281 2370
rect 1247 2246 1281 2280
rect 1247 2156 1281 2190
rect 1247 2066 1281 2100
rect 1247 1976 1281 2010
rect 1247 1886 1281 1920
rect 1247 1796 1281 1830
rect 1247 1706 1281 1740
rect 1247 1616 1281 1650
rect 1247 1526 1281 1560
rect 1247 1436 1281 1470
rect 60 1346 94 1380
rect 1247 1346 1281 1380
rect 156 1262 190 1296
rect 246 1262 280 1296
rect 336 1262 370 1296
rect 426 1262 460 1296
rect 516 1262 550 1296
rect 606 1262 640 1296
rect 696 1262 730 1296
rect 786 1262 820 1296
rect 876 1262 910 1296
rect 966 1262 1000 1296
rect 1056 1262 1090 1296
rect 1146 1262 1180 1296
rect 1402 2426 1436 2460
rect 1498 2449 1532 2483
rect 1588 2449 1622 2483
rect 1678 2449 1712 2483
rect 1768 2449 1802 2483
rect 1858 2449 1892 2483
rect 1948 2449 1982 2483
rect 2038 2449 2072 2483
rect 2128 2449 2162 2483
rect 2218 2449 2252 2483
rect 2308 2449 2342 2483
rect 2398 2449 2432 2483
rect 2488 2449 2522 2483
rect 2589 2426 2623 2460
rect 1402 2336 1436 2370
rect 1402 2246 1436 2280
rect 1402 2156 1436 2190
rect 1402 2066 1436 2100
rect 1402 1976 1436 2010
rect 1402 1886 1436 1920
rect 1402 1796 1436 1830
rect 1402 1706 1436 1740
rect 1402 1616 1436 1650
rect 1402 1526 1436 1560
rect 1402 1436 1436 1470
rect 2589 2336 2623 2370
rect 2589 2246 2623 2280
rect 2589 2156 2623 2190
rect 2589 2066 2623 2100
rect 2589 1976 2623 2010
rect 2589 1886 2623 1920
rect 2589 1796 2623 1830
rect 2589 1706 2623 1740
rect 2589 1616 2623 1650
rect 2589 1526 2623 1560
rect 2589 1436 2623 1470
rect 1402 1346 1436 1380
rect 2589 1346 2623 1380
rect 1498 1262 1532 1296
rect 1588 1262 1622 1296
rect 1678 1262 1712 1296
rect 1768 1262 1802 1296
rect 1858 1262 1892 1296
rect 1948 1262 1982 1296
rect 2038 1262 2072 1296
rect 2128 1262 2162 1296
rect 2218 1262 2252 1296
rect 2308 1262 2342 1296
rect 2398 1262 2432 1296
rect 2488 1262 2522 1296
rect 2744 2426 2778 2460
rect 2840 2449 2874 2483
rect 2930 2449 2964 2483
rect 3020 2449 3054 2483
rect 3110 2449 3144 2483
rect 3200 2449 3234 2483
rect 3290 2449 3324 2483
rect 3380 2449 3414 2483
rect 3470 2449 3504 2483
rect 3560 2449 3594 2483
rect 3650 2449 3684 2483
rect 3740 2449 3774 2483
rect 3830 2449 3864 2483
rect 3931 2426 3965 2460
rect 2744 2336 2778 2370
rect 2744 2246 2778 2280
rect 2744 2156 2778 2190
rect 2744 2066 2778 2100
rect 2744 1976 2778 2010
rect 2744 1886 2778 1920
rect 2744 1796 2778 1830
rect 2744 1706 2778 1740
rect 2744 1616 2778 1650
rect 2744 1526 2778 1560
rect 2744 1436 2778 1470
rect 3931 2336 3965 2370
rect 3931 2246 3965 2280
rect 3931 2156 3965 2190
rect 3931 2066 3965 2100
rect 3931 1976 3965 2010
rect 3931 1886 3965 1920
rect 3931 1796 3965 1830
rect 3931 1706 3965 1740
rect 3931 1616 3965 1650
rect 3931 1526 3965 1560
rect 3931 1436 3965 1470
rect 2744 1346 2778 1380
rect 3931 1346 3965 1380
rect 2840 1262 2874 1296
rect 2930 1262 2964 1296
rect 3020 1262 3054 1296
rect 3110 1262 3144 1296
rect 3200 1262 3234 1296
rect 3290 1262 3324 1296
rect 3380 1262 3414 1296
rect 3470 1262 3504 1296
rect 3560 1262 3594 1296
rect 3650 1262 3684 1296
rect 3740 1262 3774 1296
rect 3830 1262 3864 1296
rect 4086 2426 4120 2460
rect 4182 2449 4216 2483
rect 4272 2449 4306 2483
rect 4362 2449 4396 2483
rect 4452 2449 4486 2483
rect 4542 2449 4576 2483
rect 4632 2449 4666 2483
rect 4722 2449 4756 2483
rect 4812 2449 4846 2483
rect 4902 2449 4936 2483
rect 4992 2449 5026 2483
rect 5082 2449 5116 2483
rect 5172 2449 5206 2483
rect 5273 2426 5307 2460
rect 4086 2336 4120 2370
rect 4086 2246 4120 2280
rect 4086 2156 4120 2190
rect 4086 2066 4120 2100
rect 4086 1976 4120 2010
rect 4086 1886 4120 1920
rect 4086 1796 4120 1830
rect 4086 1706 4120 1740
rect 4086 1616 4120 1650
rect 4086 1526 4120 1560
rect 4086 1436 4120 1470
rect 5273 2336 5307 2370
rect 5273 2246 5307 2280
rect 5273 2156 5307 2190
rect 5273 2066 5307 2100
rect 5273 1976 5307 2010
rect 5273 1886 5307 1920
rect 5273 1796 5307 1830
rect 5273 1706 5307 1740
rect 5273 1616 5307 1650
rect 5273 1526 5307 1560
rect 5273 1436 5307 1470
rect 4086 1346 4120 1380
rect 5273 1346 5307 1380
rect 4182 1262 4216 1296
rect 4272 1262 4306 1296
rect 4362 1262 4396 1296
rect 4452 1262 4486 1296
rect 4542 1262 4576 1296
rect 4632 1262 4666 1296
rect 4722 1262 4756 1296
rect 4812 1262 4846 1296
rect 4902 1262 4936 1296
rect 4992 1262 5026 1296
rect 5082 1262 5116 1296
rect 5172 1262 5206 1296
rect 5428 2426 5462 2460
rect 5524 2449 5558 2483
rect 5614 2449 5648 2483
rect 5704 2449 5738 2483
rect 5794 2449 5828 2483
rect 5884 2449 5918 2483
rect 5974 2449 6008 2483
rect 6064 2449 6098 2483
rect 6154 2449 6188 2483
rect 6244 2449 6278 2483
rect 6334 2449 6368 2483
rect 6424 2449 6458 2483
rect 6514 2449 6548 2483
rect 6615 2426 6649 2460
rect 5428 2336 5462 2370
rect 5428 2246 5462 2280
rect 5428 2156 5462 2190
rect 5428 2066 5462 2100
rect 5428 1976 5462 2010
rect 5428 1886 5462 1920
rect 5428 1796 5462 1830
rect 5428 1706 5462 1740
rect 5428 1616 5462 1650
rect 5428 1526 5462 1560
rect 5428 1436 5462 1470
rect 6615 2336 6649 2370
rect 6615 2246 6649 2280
rect 6615 2156 6649 2190
rect 6615 2066 6649 2100
rect 6615 1976 6649 2010
rect 6615 1886 6649 1920
rect 6615 1796 6649 1830
rect 6615 1706 6649 1740
rect 6615 1616 6649 1650
rect 6615 1526 6649 1560
rect 6615 1436 6649 1470
rect 5428 1346 5462 1380
rect 6615 1346 6649 1380
rect 5524 1262 5558 1296
rect 5614 1262 5648 1296
rect 5704 1262 5738 1296
rect 5794 1262 5828 1296
rect 5884 1262 5918 1296
rect 5974 1262 6008 1296
rect 6064 1262 6098 1296
rect 6154 1262 6188 1296
rect 6244 1262 6278 1296
rect 6334 1262 6368 1296
rect 6424 1262 6458 1296
rect 6514 1262 6548 1296
rect 6770 2426 6804 2460
rect 6866 2449 6900 2483
rect 6956 2449 6990 2483
rect 7046 2449 7080 2483
rect 7136 2449 7170 2483
rect 7226 2449 7260 2483
rect 7316 2449 7350 2483
rect 7406 2449 7440 2483
rect 7496 2449 7530 2483
rect 7586 2449 7620 2483
rect 7676 2449 7710 2483
rect 7766 2449 7800 2483
rect 7856 2449 7890 2483
rect 7957 2426 7991 2460
rect 6770 2336 6804 2370
rect 6770 2246 6804 2280
rect 6770 2156 6804 2190
rect 6770 2066 6804 2100
rect 6770 1976 6804 2010
rect 6770 1886 6804 1920
rect 6770 1796 6804 1830
rect 6770 1706 6804 1740
rect 6770 1616 6804 1650
rect 6770 1526 6804 1560
rect 6770 1436 6804 1470
rect 7957 2336 7991 2370
rect 7957 2246 7991 2280
rect 7957 2156 7991 2190
rect 7957 2066 7991 2100
rect 7957 1976 7991 2010
rect 7957 1886 7991 1920
rect 7957 1796 7991 1830
rect 7957 1706 7991 1740
rect 7957 1616 7991 1650
rect 7957 1526 7991 1560
rect 7957 1436 7991 1470
rect 6770 1346 6804 1380
rect 7957 1346 7991 1380
rect 6866 1262 6900 1296
rect 6956 1262 6990 1296
rect 7046 1262 7080 1296
rect 7136 1262 7170 1296
rect 7226 1262 7260 1296
rect 7316 1262 7350 1296
rect 7406 1262 7440 1296
rect 7496 1262 7530 1296
rect 7586 1262 7620 1296
rect 7676 1262 7710 1296
rect 7766 1262 7800 1296
rect 7856 1262 7890 1296
rect 8112 2426 8146 2460
rect 8208 2449 8242 2483
rect 8298 2449 8332 2483
rect 8388 2449 8422 2483
rect 8478 2449 8512 2483
rect 8568 2449 8602 2483
rect 8658 2449 8692 2483
rect 8748 2449 8782 2483
rect 8838 2449 8872 2483
rect 8928 2449 8962 2483
rect 9018 2449 9052 2483
rect 9108 2449 9142 2483
rect 9198 2449 9232 2483
rect 9299 2426 9333 2460
rect 8112 2336 8146 2370
rect 8112 2246 8146 2280
rect 8112 2156 8146 2190
rect 8112 2066 8146 2100
rect 8112 1976 8146 2010
rect 8112 1886 8146 1920
rect 8112 1796 8146 1830
rect 8112 1706 8146 1740
rect 8112 1616 8146 1650
rect 8112 1526 8146 1560
rect 8112 1436 8146 1470
rect 9299 2336 9333 2370
rect 9299 2246 9333 2280
rect 9299 2156 9333 2190
rect 9299 2066 9333 2100
rect 9299 1976 9333 2010
rect 9299 1886 9333 1920
rect 9299 1796 9333 1830
rect 9299 1706 9333 1740
rect 9299 1616 9333 1650
rect 9299 1526 9333 1560
rect 9299 1436 9333 1470
rect 8112 1346 8146 1380
rect 9299 1346 9333 1380
rect 8208 1262 8242 1296
rect 8298 1262 8332 1296
rect 8388 1262 8422 1296
rect 8478 1262 8512 1296
rect 8568 1262 8602 1296
rect 8658 1262 8692 1296
rect 8748 1262 8782 1296
rect 8838 1262 8872 1296
rect 8928 1262 8962 1296
rect 9018 1262 9052 1296
rect 9108 1262 9142 1296
rect 9198 1262 9232 1296
rect 6770 1084 6804 1118
rect 6866 1107 6900 1141
rect 6956 1107 6990 1141
rect 7046 1107 7080 1141
rect 7136 1107 7170 1141
rect 7226 1107 7260 1141
rect 7316 1107 7350 1141
rect 7406 1107 7440 1141
rect 7496 1107 7530 1141
rect 7586 1107 7620 1141
rect 7676 1107 7710 1141
rect 7766 1107 7800 1141
rect 7856 1107 7890 1141
rect 7957 1084 7991 1118
rect 6770 994 6804 1028
rect 6770 904 6804 938
rect 6770 814 6804 848
rect 6770 724 6804 758
rect 6770 634 6804 668
rect 6770 544 6804 578
rect 6770 454 6804 488
rect 6770 364 6804 398
rect 6770 274 6804 308
rect 6770 184 6804 218
rect 6770 94 6804 128
rect 7957 994 7991 1028
rect 7957 904 7991 938
rect 7957 814 7991 848
rect 7957 724 7991 758
rect 7957 634 7991 668
rect 7957 544 7991 578
rect 7957 454 7991 488
rect 7957 364 7991 398
rect 7957 274 7991 308
rect 7957 184 7991 218
rect 7957 94 7991 128
rect 6770 4 6804 38
rect 7957 4 7991 38
rect 6866 -80 6900 -46
rect 6956 -80 6990 -46
rect 7046 -80 7080 -46
rect 7136 -80 7170 -46
rect 7226 -80 7260 -46
rect 7316 -80 7350 -46
rect 7406 -80 7440 -46
rect 7496 -80 7530 -46
rect 7586 -80 7620 -46
rect 7676 -80 7710 -46
rect 7766 -80 7800 -46
rect 7856 -80 7890 -46
rect 8112 1084 8146 1118
rect 8208 1107 8242 1141
rect 8298 1107 8332 1141
rect 8388 1107 8422 1141
rect 8478 1107 8512 1141
rect 8568 1107 8602 1141
rect 8658 1107 8692 1141
rect 8748 1107 8782 1141
rect 8838 1107 8872 1141
rect 8928 1107 8962 1141
rect 9018 1107 9052 1141
rect 9108 1107 9142 1141
rect 9198 1107 9232 1141
rect 9299 1084 9333 1118
rect 8112 994 8146 1028
rect 8112 904 8146 938
rect 8112 814 8146 848
rect 8112 724 8146 758
rect 8112 634 8146 668
rect 8112 544 8146 578
rect 8112 454 8146 488
rect 8112 364 8146 398
rect 8112 274 8146 308
rect 8112 184 8146 218
rect 8112 94 8146 128
rect 9299 994 9333 1028
rect 9299 904 9333 938
rect 9299 814 9333 848
rect 9299 724 9333 758
rect 9299 634 9333 668
rect 9299 544 9333 578
rect 9299 454 9333 488
rect 9299 364 9333 398
rect 9299 274 9333 308
rect 9299 184 9333 218
rect 9299 94 9333 128
rect 8112 4 8146 38
rect 9299 4 9333 38
rect 8208 -80 8242 -46
rect 8298 -80 8332 -46
rect 8388 -80 8422 -46
rect 8478 -80 8512 -46
rect 8568 -80 8602 -46
rect 8658 -80 8692 -46
rect 8748 -80 8782 -46
rect 8838 -80 8872 -46
rect 8928 -80 8962 -46
rect 9018 -80 9052 -46
rect 9108 -80 9142 -46
rect 9198 -80 9232 -46
rect 6770 -258 6804 -224
rect 6866 -235 6900 -201
rect 6956 -235 6990 -201
rect 7046 -235 7080 -201
rect 7136 -235 7170 -201
rect 7226 -235 7260 -201
rect 7316 -235 7350 -201
rect 7406 -235 7440 -201
rect 7496 -235 7530 -201
rect 7586 -235 7620 -201
rect 7676 -235 7710 -201
rect 7766 -235 7800 -201
rect 7856 -235 7890 -201
rect 7957 -258 7991 -224
rect 6770 -348 6804 -314
rect 6770 -438 6804 -404
rect 6770 -528 6804 -494
rect 6770 -618 6804 -584
rect 6770 -708 6804 -674
rect 6770 -798 6804 -764
rect 6770 -888 6804 -854
rect 6770 -978 6804 -944
rect 6770 -1068 6804 -1034
rect 6770 -1158 6804 -1124
rect 6770 -1248 6804 -1214
rect 7957 -348 7991 -314
rect 7957 -438 7991 -404
rect 7957 -528 7991 -494
rect 7957 -618 7991 -584
rect 7957 -708 7991 -674
rect 7957 -798 7991 -764
rect 7957 -888 7991 -854
rect 7957 -978 7991 -944
rect 7957 -1068 7991 -1034
rect 7957 -1158 7991 -1124
rect 7957 -1248 7991 -1214
rect 6770 -1338 6804 -1304
rect 7957 -1338 7991 -1304
rect 6866 -1422 6900 -1388
rect 6956 -1422 6990 -1388
rect 7046 -1422 7080 -1388
rect 7136 -1422 7170 -1388
rect 7226 -1422 7260 -1388
rect 7316 -1422 7350 -1388
rect 7406 -1422 7440 -1388
rect 7496 -1422 7530 -1388
rect 7586 -1422 7620 -1388
rect 7676 -1422 7710 -1388
rect 7766 -1422 7800 -1388
rect 7856 -1422 7890 -1388
rect 8112 -258 8146 -224
rect 8208 -235 8242 -201
rect 8298 -235 8332 -201
rect 8388 -235 8422 -201
rect 8478 -235 8512 -201
rect 8568 -235 8602 -201
rect 8658 -235 8692 -201
rect 8748 -235 8782 -201
rect 8838 -235 8872 -201
rect 8928 -235 8962 -201
rect 9018 -235 9052 -201
rect 9108 -235 9142 -201
rect 9198 -235 9232 -201
rect 9299 -258 9333 -224
rect 8112 -348 8146 -314
rect 8112 -438 8146 -404
rect 8112 -528 8146 -494
rect 8112 -618 8146 -584
rect 8112 -708 8146 -674
rect 8112 -798 8146 -764
rect 8112 -888 8146 -854
rect 8112 -978 8146 -944
rect 8112 -1068 8146 -1034
rect 8112 -1158 8146 -1124
rect 8112 -1248 8146 -1214
rect 9299 -348 9333 -314
rect 9299 -438 9333 -404
rect 9299 -528 9333 -494
rect 9299 -618 9333 -584
rect 9299 -708 9333 -674
rect 9299 -798 9333 -764
rect 9299 -888 9333 -854
rect 9299 -978 9333 -944
rect 9299 -1068 9333 -1034
rect 9299 -1158 9333 -1124
rect 9299 -1248 9333 -1214
rect 8112 -1338 8146 -1304
rect 9299 -1338 9333 -1304
rect 8208 -1422 8242 -1388
rect 8298 -1422 8332 -1388
rect 8388 -1422 8422 -1388
rect 8478 -1422 8512 -1388
rect 8568 -1422 8602 -1388
rect 8658 -1422 8692 -1388
rect 8748 -1422 8782 -1388
rect 8838 -1422 8872 -1388
rect 8928 -1422 8962 -1388
rect 9018 -1422 9052 -1388
rect 9108 -1422 9142 -1388
rect 9198 -1422 9232 -1388
<< nsubdiffcont >>
rect 320 3644 354 3678
rect 410 3644 444 3678
rect 500 3644 534 3678
rect 590 3644 624 3678
rect 680 3644 714 3678
rect 770 3644 804 3678
rect 860 3644 894 3678
rect 950 3644 984 3678
rect 1040 3644 1074 3678
rect 208 3587 242 3621
rect 1098 3568 1132 3602
rect 208 3497 242 3531
rect 208 3407 242 3441
rect 208 3317 242 3351
rect 208 3227 242 3261
rect 208 3137 242 3171
rect 208 3047 242 3081
rect 208 2957 242 2991
rect 208 2867 242 2901
rect 1098 3478 1132 3512
rect 1098 3388 1132 3422
rect 1098 3298 1132 3332
rect 1098 3208 1132 3242
rect 1098 3118 1132 3152
rect 1098 3028 1132 3062
rect 1098 2938 1132 2972
rect 1098 2848 1132 2882
rect 286 2754 320 2788
rect 376 2754 410 2788
rect 466 2754 500 2788
rect 556 2754 590 2788
rect 646 2754 680 2788
rect 736 2754 770 2788
rect 826 2754 860 2788
rect 916 2754 950 2788
rect 1006 2754 1040 2788
rect 1662 3644 1696 3678
rect 1752 3644 1786 3678
rect 1842 3644 1876 3678
rect 1932 3644 1966 3678
rect 2022 3644 2056 3678
rect 2112 3644 2146 3678
rect 2202 3644 2236 3678
rect 2292 3644 2326 3678
rect 2382 3644 2416 3678
rect 1550 3587 1584 3621
rect 2440 3568 2474 3602
rect 1550 3497 1584 3531
rect 1550 3407 1584 3441
rect 1550 3317 1584 3351
rect 1550 3227 1584 3261
rect 1550 3137 1584 3171
rect 1550 3047 1584 3081
rect 1550 2957 1584 2991
rect 1550 2867 1584 2901
rect 2440 3478 2474 3512
rect 2440 3388 2474 3422
rect 2440 3298 2474 3332
rect 2440 3208 2474 3242
rect 2440 3118 2474 3152
rect 2440 3028 2474 3062
rect 2440 2938 2474 2972
rect 2440 2848 2474 2882
rect 1628 2754 1662 2788
rect 1718 2754 1752 2788
rect 1808 2754 1842 2788
rect 1898 2754 1932 2788
rect 1988 2754 2022 2788
rect 2078 2754 2112 2788
rect 2168 2754 2202 2788
rect 2258 2754 2292 2788
rect 2348 2754 2382 2788
rect 3004 3644 3038 3678
rect 3094 3644 3128 3678
rect 3184 3644 3218 3678
rect 3274 3644 3308 3678
rect 3364 3644 3398 3678
rect 3454 3644 3488 3678
rect 3544 3644 3578 3678
rect 3634 3644 3668 3678
rect 3724 3644 3758 3678
rect 2892 3587 2926 3621
rect 3782 3568 3816 3602
rect 2892 3497 2926 3531
rect 2892 3407 2926 3441
rect 2892 3317 2926 3351
rect 2892 3227 2926 3261
rect 2892 3137 2926 3171
rect 2892 3047 2926 3081
rect 2892 2957 2926 2991
rect 2892 2867 2926 2901
rect 3782 3478 3816 3512
rect 3782 3388 3816 3422
rect 3782 3298 3816 3332
rect 3782 3208 3816 3242
rect 3782 3118 3816 3152
rect 3782 3028 3816 3062
rect 3782 2938 3816 2972
rect 3782 2848 3816 2882
rect 2970 2754 3004 2788
rect 3060 2754 3094 2788
rect 3150 2754 3184 2788
rect 3240 2754 3274 2788
rect 3330 2754 3364 2788
rect 3420 2754 3454 2788
rect 3510 2754 3544 2788
rect 3600 2754 3634 2788
rect 3690 2754 3724 2788
rect 4346 3644 4380 3678
rect 4436 3644 4470 3678
rect 4526 3644 4560 3678
rect 4616 3644 4650 3678
rect 4706 3644 4740 3678
rect 4796 3644 4830 3678
rect 4886 3644 4920 3678
rect 4976 3644 5010 3678
rect 5066 3644 5100 3678
rect 4234 3587 4268 3621
rect 5124 3568 5158 3602
rect 4234 3497 4268 3531
rect 4234 3407 4268 3441
rect 4234 3317 4268 3351
rect 4234 3227 4268 3261
rect 4234 3137 4268 3171
rect 4234 3047 4268 3081
rect 4234 2957 4268 2991
rect 4234 2867 4268 2901
rect 5124 3478 5158 3512
rect 5124 3388 5158 3422
rect 5124 3298 5158 3332
rect 5124 3208 5158 3242
rect 5124 3118 5158 3152
rect 5124 3028 5158 3062
rect 5124 2938 5158 2972
rect 5124 2848 5158 2882
rect 4312 2754 4346 2788
rect 4402 2754 4436 2788
rect 4492 2754 4526 2788
rect 4582 2754 4616 2788
rect 4672 2754 4706 2788
rect 4762 2754 4796 2788
rect 4852 2754 4886 2788
rect 4942 2754 4976 2788
rect 5032 2754 5066 2788
rect 5688 3644 5722 3678
rect 5778 3644 5812 3678
rect 5868 3644 5902 3678
rect 5958 3644 5992 3678
rect 6048 3644 6082 3678
rect 6138 3644 6172 3678
rect 6228 3644 6262 3678
rect 6318 3644 6352 3678
rect 6408 3644 6442 3678
rect 5576 3587 5610 3621
rect 6466 3568 6500 3602
rect 5576 3497 5610 3531
rect 5576 3407 5610 3441
rect 5576 3317 5610 3351
rect 5576 3227 5610 3261
rect 5576 3137 5610 3171
rect 5576 3047 5610 3081
rect 5576 2957 5610 2991
rect 5576 2867 5610 2901
rect 6466 3478 6500 3512
rect 6466 3388 6500 3422
rect 6466 3298 6500 3332
rect 6466 3208 6500 3242
rect 6466 3118 6500 3152
rect 6466 3028 6500 3062
rect 6466 2938 6500 2972
rect 6466 2848 6500 2882
rect 5654 2754 5688 2788
rect 5744 2754 5778 2788
rect 5834 2754 5868 2788
rect 5924 2754 5958 2788
rect 6014 2754 6048 2788
rect 6104 2754 6138 2788
rect 6194 2754 6228 2788
rect 6284 2754 6318 2788
rect 6374 2754 6408 2788
rect 7030 3644 7064 3678
rect 7120 3644 7154 3678
rect 7210 3644 7244 3678
rect 7300 3644 7334 3678
rect 7390 3644 7424 3678
rect 7480 3644 7514 3678
rect 7570 3644 7604 3678
rect 7660 3644 7694 3678
rect 7750 3644 7784 3678
rect 6918 3587 6952 3621
rect 7808 3568 7842 3602
rect 6918 3497 6952 3531
rect 6918 3407 6952 3441
rect 6918 3317 6952 3351
rect 6918 3227 6952 3261
rect 6918 3137 6952 3171
rect 6918 3047 6952 3081
rect 6918 2957 6952 2991
rect 6918 2867 6952 2901
rect 7808 3478 7842 3512
rect 7808 3388 7842 3422
rect 7808 3298 7842 3332
rect 7808 3208 7842 3242
rect 7808 3118 7842 3152
rect 7808 3028 7842 3062
rect 7808 2938 7842 2972
rect 7808 2848 7842 2882
rect 6996 2754 7030 2788
rect 7086 2754 7120 2788
rect 7176 2754 7210 2788
rect 7266 2754 7300 2788
rect 7356 2754 7390 2788
rect 7446 2754 7480 2788
rect 7536 2754 7570 2788
rect 7626 2754 7660 2788
rect 7716 2754 7750 2788
rect 8372 3644 8406 3678
rect 8462 3644 8496 3678
rect 8552 3644 8586 3678
rect 8642 3644 8676 3678
rect 8732 3644 8766 3678
rect 8822 3644 8856 3678
rect 8912 3644 8946 3678
rect 9002 3644 9036 3678
rect 9092 3644 9126 3678
rect 8260 3587 8294 3621
rect 9150 3568 9184 3602
rect 8260 3497 8294 3531
rect 8260 3407 8294 3441
rect 8260 3317 8294 3351
rect 8260 3227 8294 3261
rect 8260 3137 8294 3171
rect 8260 3047 8294 3081
rect 8260 2957 8294 2991
rect 8260 2867 8294 2901
rect 9150 3478 9184 3512
rect 9150 3388 9184 3422
rect 9150 3298 9184 3332
rect 9150 3208 9184 3242
rect 9150 3118 9184 3152
rect 9150 3028 9184 3062
rect 9150 2938 9184 2972
rect 9150 2848 9184 2882
rect 8338 2754 8372 2788
rect 8428 2754 8462 2788
rect 8518 2754 8552 2788
rect 8608 2754 8642 2788
rect 8698 2754 8732 2788
rect 8788 2754 8822 2788
rect 8878 2754 8912 2788
rect 8968 2754 9002 2788
rect 9058 2754 9092 2788
rect 320 2302 354 2336
rect 410 2302 444 2336
rect 500 2302 534 2336
rect 590 2302 624 2336
rect 680 2302 714 2336
rect 770 2302 804 2336
rect 860 2302 894 2336
rect 950 2302 984 2336
rect 1040 2302 1074 2336
rect 208 2245 242 2279
rect 1098 2226 1132 2260
rect 208 2155 242 2189
rect 208 2065 242 2099
rect 208 1975 242 2009
rect 208 1885 242 1919
rect 208 1795 242 1829
rect 208 1705 242 1739
rect 208 1615 242 1649
rect 208 1525 242 1559
rect 1098 2136 1132 2170
rect 1098 2046 1132 2080
rect 1098 1956 1132 1990
rect 1098 1866 1132 1900
rect 1098 1776 1132 1810
rect 1098 1686 1132 1720
rect 1098 1596 1132 1630
rect 1098 1506 1132 1540
rect 286 1412 320 1446
rect 376 1412 410 1446
rect 466 1412 500 1446
rect 556 1412 590 1446
rect 646 1412 680 1446
rect 736 1412 770 1446
rect 826 1412 860 1446
rect 916 1412 950 1446
rect 1006 1412 1040 1446
rect 1662 2302 1696 2336
rect 1752 2302 1786 2336
rect 1842 2302 1876 2336
rect 1932 2302 1966 2336
rect 2022 2302 2056 2336
rect 2112 2302 2146 2336
rect 2202 2302 2236 2336
rect 2292 2302 2326 2336
rect 2382 2302 2416 2336
rect 1550 2245 1584 2279
rect 2440 2226 2474 2260
rect 1550 2155 1584 2189
rect 1550 2065 1584 2099
rect 1550 1975 1584 2009
rect 1550 1885 1584 1919
rect 1550 1795 1584 1829
rect 1550 1705 1584 1739
rect 1550 1615 1584 1649
rect 1550 1525 1584 1559
rect 2440 2136 2474 2170
rect 2440 2046 2474 2080
rect 2440 1956 2474 1990
rect 2440 1866 2474 1900
rect 2440 1776 2474 1810
rect 2440 1686 2474 1720
rect 2440 1596 2474 1630
rect 2440 1506 2474 1540
rect 1628 1412 1662 1446
rect 1718 1412 1752 1446
rect 1808 1412 1842 1446
rect 1898 1412 1932 1446
rect 1988 1412 2022 1446
rect 2078 1412 2112 1446
rect 2168 1412 2202 1446
rect 2258 1412 2292 1446
rect 2348 1412 2382 1446
rect 3004 2302 3038 2336
rect 3094 2302 3128 2336
rect 3184 2302 3218 2336
rect 3274 2302 3308 2336
rect 3364 2302 3398 2336
rect 3454 2302 3488 2336
rect 3544 2302 3578 2336
rect 3634 2302 3668 2336
rect 3724 2302 3758 2336
rect 2892 2245 2926 2279
rect 3782 2226 3816 2260
rect 2892 2155 2926 2189
rect 2892 2065 2926 2099
rect 2892 1975 2926 2009
rect 2892 1885 2926 1919
rect 2892 1795 2926 1829
rect 2892 1705 2926 1739
rect 2892 1615 2926 1649
rect 2892 1525 2926 1559
rect 3782 2136 3816 2170
rect 3782 2046 3816 2080
rect 3782 1956 3816 1990
rect 3782 1866 3816 1900
rect 3782 1776 3816 1810
rect 3782 1686 3816 1720
rect 3782 1596 3816 1630
rect 3782 1506 3816 1540
rect 2970 1412 3004 1446
rect 3060 1412 3094 1446
rect 3150 1412 3184 1446
rect 3240 1412 3274 1446
rect 3330 1412 3364 1446
rect 3420 1412 3454 1446
rect 3510 1412 3544 1446
rect 3600 1412 3634 1446
rect 3690 1412 3724 1446
rect 4346 2302 4380 2336
rect 4436 2302 4470 2336
rect 4526 2302 4560 2336
rect 4616 2302 4650 2336
rect 4706 2302 4740 2336
rect 4796 2302 4830 2336
rect 4886 2302 4920 2336
rect 4976 2302 5010 2336
rect 5066 2302 5100 2336
rect 4234 2245 4268 2279
rect 5124 2226 5158 2260
rect 4234 2155 4268 2189
rect 4234 2065 4268 2099
rect 4234 1975 4268 2009
rect 4234 1885 4268 1919
rect 4234 1795 4268 1829
rect 4234 1705 4268 1739
rect 4234 1615 4268 1649
rect 4234 1525 4268 1559
rect 5124 2136 5158 2170
rect 5124 2046 5158 2080
rect 5124 1956 5158 1990
rect 5124 1866 5158 1900
rect 5124 1776 5158 1810
rect 5124 1686 5158 1720
rect 5124 1596 5158 1630
rect 5124 1506 5158 1540
rect 4312 1412 4346 1446
rect 4402 1412 4436 1446
rect 4492 1412 4526 1446
rect 4582 1412 4616 1446
rect 4672 1412 4706 1446
rect 4762 1412 4796 1446
rect 4852 1412 4886 1446
rect 4942 1412 4976 1446
rect 5032 1412 5066 1446
rect 5688 2302 5722 2336
rect 5778 2302 5812 2336
rect 5868 2302 5902 2336
rect 5958 2302 5992 2336
rect 6048 2302 6082 2336
rect 6138 2302 6172 2336
rect 6228 2302 6262 2336
rect 6318 2302 6352 2336
rect 6408 2302 6442 2336
rect 5576 2245 5610 2279
rect 6466 2226 6500 2260
rect 5576 2155 5610 2189
rect 5576 2065 5610 2099
rect 5576 1975 5610 2009
rect 5576 1885 5610 1919
rect 5576 1795 5610 1829
rect 5576 1705 5610 1739
rect 5576 1615 5610 1649
rect 5576 1525 5610 1559
rect 6466 2136 6500 2170
rect 6466 2046 6500 2080
rect 6466 1956 6500 1990
rect 6466 1866 6500 1900
rect 6466 1776 6500 1810
rect 6466 1686 6500 1720
rect 6466 1596 6500 1630
rect 6466 1506 6500 1540
rect 5654 1412 5688 1446
rect 5744 1412 5778 1446
rect 5834 1412 5868 1446
rect 5924 1412 5958 1446
rect 6014 1412 6048 1446
rect 6104 1412 6138 1446
rect 6194 1412 6228 1446
rect 6284 1412 6318 1446
rect 6374 1412 6408 1446
rect 7030 2302 7064 2336
rect 7120 2302 7154 2336
rect 7210 2302 7244 2336
rect 7300 2302 7334 2336
rect 7390 2302 7424 2336
rect 7480 2302 7514 2336
rect 7570 2302 7604 2336
rect 7660 2302 7694 2336
rect 7750 2302 7784 2336
rect 6918 2245 6952 2279
rect 7808 2226 7842 2260
rect 6918 2155 6952 2189
rect 6918 2065 6952 2099
rect 6918 1975 6952 2009
rect 6918 1885 6952 1919
rect 6918 1795 6952 1829
rect 6918 1705 6952 1739
rect 6918 1615 6952 1649
rect 6918 1525 6952 1559
rect 7808 2136 7842 2170
rect 7808 2046 7842 2080
rect 7808 1956 7842 1990
rect 7808 1866 7842 1900
rect 7808 1776 7842 1810
rect 7808 1686 7842 1720
rect 7808 1596 7842 1630
rect 7808 1506 7842 1540
rect 6996 1412 7030 1446
rect 7086 1412 7120 1446
rect 7176 1412 7210 1446
rect 7266 1412 7300 1446
rect 7356 1412 7390 1446
rect 7446 1412 7480 1446
rect 7536 1412 7570 1446
rect 7626 1412 7660 1446
rect 7716 1412 7750 1446
rect 8372 2302 8406 2336
rect 8462 2302 8496 2336
rect 8552 2302 8586 2336
rect 8642 2302 8676 2336
rect 8732 2302 8766 2336
rect 8822 2302 8856 2336
rect 8912 2302 8946 2336
rect 9002 2302 9036 2336
rect 9092 2302 9126 2336
rect 8260 2245 8294 2279
rect 9150 2226 9184 2260
rect 8260 2155 8294 2189
rect 8260 2065 8294 2099
rect 8260 1975 8294 2009
rect 8260 1885 8294 1919
rect 8260 1795 8294 1829
rect 8260 1705 8294 1739
rect 8260 1615 8294 1649
rect 8260 1525 8294 1559
rect 9150 2136 9184 2170
rect 9150 2046 9184 2080
rect 9150 1956 9184 1990
rect 9150 1866 9184 1900
rect 9150 1776 9184 1810
rect 9150 1686 9184 1720
rect 9150 1596 9184 1630
rect 9150 1506 9184 1540
rect 8338 1412 8372 1446
rect 8428 1412 8462 1446
rect 8518 1412 8552 1446
rect 8608 1412 8642 1446
rect 8698 1412 8732 1446
rect 8788 1412 8822 1446
rect 8878 1412 8912 1446
rect 8968 1412 9002 1446
rect 9058 1412 9092 1446
rect 7030 960 7064 994
rect 7120 960 7154 994
rect 7210 960 7244 994
rect 7300 960 7334 994
rect 7390 960 7424 994
rect 7480 960 7514 994
rect 7570 960 7604 994
rect 7660 960 7694 994
rect 7750 960 7784 994
rect 6918 903 6952 937
rect 7808 884 7842 918
rect 6918 813 6952 847
rect 6918 723 6952 757
rect 6918 633 6952 667
rect 6918 543 6952 577
rect 6918 453 6952 487
rect 6918 363 6952 397
rect 6918 273 6952 307
rect 6918 183 6952 217
rect 7808 794 7842 828
rect 7808 704 7842 738
rect 7808 614 7842 648
rect 7808 524 7842 558
rect 7808 434 7842 468
rect 7808 344 7842 378
rect 7808 254 7842 288
rect 7808 164 7842 198
rect 6996 70 7030 104
rect 7086 70 7120 104
rect 7176 70 7210 104
rect 7266 70 7300 104
rect 7356 70 7390 104
rect 7446 70 7480 104
rect 7536 70 7570 104
rect 7626 70 7660 104
rect 7716 70 7750 104
rect 8372 960 8406 994
rect 8462 960 8496 994
rect 8552 960 8586 994
rect 8642 960 8676 994
rect 8732 960 8766 994
rect 8822 960 8856 994
rect 8912 960 8946 994
rect 9002 960 9036 994
rect 9092 960 9126 994
rect 8260 903 8294 937
rect 9150 884 9184 918
rect 8260 813 8294 847
rect 8260 723 8294 757
rect 8260 633 8294 667
rect 8260 543 8294 577
rect 8260 453 8294 487
rect 8260 363 8294 397
rect 8260 273 8294 307
rect 8260 183 8294 217
rect 9150 794 9184 828
rect 9150 704 9184 738
rect 9150 614 9184 648
rect 9150 524 9184 558
rect 9150 434 9184 468
rect 9150 344 9184 378
rect 9150 254 9184 288
rect 9150 164 9184 198
rect 8338 70 8372 104
rect 8428 70 8462 104
rect 8518 70 8552 104
rect 8608 70 8642 104
rect 8698 70 8732 104
rect 8788 70 8822 104
rect 8878 70 8912 104
rect 8968 70 9002 104
rect 9058 70 9092 104
rect 7030 -382 7064 -348
rect 7120 -382 7154 -348
rect 7210 -382 7244 -348
rect 7300 -382 7334 -348
rect 7390 -382 7424 -348
rect 7480 -382 7514 -348
rect 7570 -382 7604 -348
rect 7660 -382 7694 -348
rect 7750 -382 7784 -348
rect 6918 -439 6952 -405
rect 7808 -458 7842 -424
rect 6918 -529 6952 -495
rect 6918 -619 6952 -585
rect 6918 -709 6952 -675
rect 6918 -799 6952 -765
rect 6918 -889 6952 -855
rect 6918 -979 6952 -945
rect 6918 -1069 6952 -1035
rect 6918 -1159 6952 -1125
rect 7808 -548 7842 -514
rect 7808 -638 7842 -604
rect 7808 -728 7842 -694
rect 7808 -818 7842 -784
rect 7808 -908 7842 -874
rect 7808 -998 7842 -964
rect 7808 -1088 7842 -1054
rect 7808 -1178 7842 -1144
rect 6996 -1272 7030 -1238
rect 7086 -1272 7120 -1238
rect 7176 -1272 7210 -1238
rect 7266 -1272 7300 -1238
rect 7356 -1272 7390 -1238
rect 7446 -1272 7480 -1238
rect 7536 -1272 7570 -1238
rect 7626 -1272 7660 -1238
rect 7716 -1272 7750 -1238
rect 8372 -382 8406 -348
rect 8462 -382 8496 -348
rect 8552 -382 8586 -348
rect 8642 -382 8676 -348
rect 8732 -382 8766 -348
rect 8822 -382 8856 -348
rect 8912 -382 8946 -348
rect 9002 -382 9036 -348
rect 9092 -382 9126 -348
rect 8260 -439 8294 -405
rect 9150 -458 9184 -424
rect 8260 -529 8294 -495
rect 8260 -619 8294 -585
rect 8260 -709 8294 -675
rect 8260 -799 8294 -765
rect 8260 -889 8294 -855
rect 8260 -979 8294 -945
rect 8260 -1069 8294 -1035
rect 8260 -1159 8294 -1125
rect 9150 -548 9184 -514
rect 9150 -638 9184 -604
rect 9150 -728 9184 -694
rect 9150 -818 9184 -784
rect 9150 -908 9184 -874
rect 9150 -998 9184 -964
rect 9150 -1088 9184 -1054
rect 9150 -1178 9184 -1144
rect 8338 -1272 8372 -1238
rect 8428 -1272 8462 -1238
rect 8518 -1272 8552 -1238
rect 8608 -1272 8642 -1238
rect 8698 -1272 8732 -1238
rect 8788 -1272 8822 -1238
rect 8878 -1272 8912 -1238
rect 8968 -1272 9002 -1238
rect 9058 -1272 9092 -1238
<< locali >>
rect 1112 3860 1525 3864
rect 26 3850 334 3860
rect 1112 3850 9366 3860
rect 26 3838 9366 3850
rect 26 3825 379 3838
rect 965 3825 9366 3838
rect 26 3802 156 3825
rect 26 3768 60 3802
rect 94 3791 156 3802
rect 190 3791 246 3825
rect 280 3791 336 3825
rect 370 3791 379 3825
rect 965 3791 966 3825
rect 1000 3791 1056 3825
rect 1090 3791 1146 3825
rect 1180 3802 1498 3825
rect 1180 3791 1247 3802
rect 94 3768 379 3791
rect 26 3712 379 3768
rect 26 3678 60 3712
rect 94 3678 379 3712
rect 965 3768 1247 3791
rect 1281 3768 1402 3802
rect 1436 3791 1498 3802
rect 1532 3791 1588 3825
rect 1622 3791 1678 3825
rect 1712 3791 1768 3825
rect 1802 3791 1858 3825
rect 1892 3791 1948 3825
rect 1982 3791 2038 3825
rect 2072 3791 2128 3825
rect 2162 3791 2218 3825
rect 2252 3791 2308 3825
rect 2342 3791 2398 3825
rect 2432 3791 2488 3825
rect 2522 3802 2840 3825
rect 2522 3791 2589 3802
rect 1436 3768 2589 3791
rect 2623 3768 2744 3802
rect 2778 3791 2840 3802
rect 2874 3791 2930 3825
rect 2964 3791 3020 3825
rect 3054 3791 3110 3825
rect 3144 3791 3200 3825
rect 3234 3791 3290 3825
rect 3324 3791 3380 3825
rect 3414 3791 3470 3825
rect 3504 3791 3560 3825
rect 3594 3791 3650 3825
rect 3684 3791 3740 3825
rect 3774 3791 3830 3825
rect 3864 3802 4182 3825
rect 3864 3791 3931 3802
rect 2778 3768 3931 3791
rect 3965 3768 4086 3802
rect 4120 3791 4182 3802
rect 4216 3791 4272 3825
rect 4306 3791 4362 3825
rect 4396 3791 4452 3825
rect 4486 3791 4542 3825
rect 4576 3791 4632 3825
rect 4666 3791 4722 3825
rect 4756 3791 4812 3825
rect 4846 3791 4902 3825
rect 4936 3791 4992 3825
rect 5026 3791 5082 3825
rect 5116 3791 5172 3825
rect 5206 3802 5524 3825
rect 5206 3791 5273 3802
rect 4120 3768 5273 3791
rect 5307 3768 5428 3802
rect 5462 3791 5524 3802
rect 5558 3791 5614 3825
rect 5648 3791 5704 3825
rect 5738 3791 5794 3825
rect 5828 3791 5884 3825
rect 5918 3791 5974 3825
rect 6008 3791 6064 3825
rect 6098 3791 6154 3825
rect 6188 3791 6244 3825
rect 6278 3791 6334 3825
rect 6368 3791 6424 3825
rect 6458 3791 6514 3825
rect 6548 3802 6866 3825
rect 6548 3791 6615 3802
rect 5462 3768 6615 3791
rect 6649 3768 6770 3802
rect 6804 3791 6866 3802
rect 6900 3791 6956 3825
rect 6990 3791 7046 3825
rect 7080 3791 7136 3825
rect 7170 3791 7226 3825
rect 7260 3791 7316 3825
rect 7350 3791 7406 3825
rect 7440 3791 7496 3825
rect 7530 3791 7586 3825
rect 7620 3791 7676 3825
rect 7710 3791 7766 3825
rect 7800 3791 7856 3825
rect 7890 3802 8208 3825
rect 7890 3791 7957 3802
rect 6804 3768 7957 3791
rect 7991 3768 8112 3802
rect 8146 3791 8208 3802
rect 8242 3791 8298 3825
rect 8332 3791 8388 3825
rect 8422 3791 8478 3825
rect 8512 3791 8568 3825
rect 8602 3791 8658 3825
rect 8692 3791 8748 3825
rect 8782 3791 8838 3825
rect 8872 3791 8928 3825
rect 8962 3791 9018 3825
rect 9052 3791 9108 3825
rect 9142 3791 9198 3825
rect 9232 3802 9366 3825
rect 9232 3791 9299 3802
rect 8146 3768 9299 3791
rect 9333 3768 9366 3802
rect 965 3712 9366 3768
rect 965 3678 1247 3712
rect 1281 3678 1402 3712
rect 1436 3678 2589 3712
rect 2623 3678 2744 3712
rect 2778 3678 3931 3712
rect 3965 3678 4086 3712
rect 4120 3678 5273 3712
rect 5307 3678 5428 3712
rect 5462 3678 6615 3712
rect 6649 3678 6770 3712
rect 6804 3678 7957 3712
rect 7991 3678 8112 3712
rect 8146 3678 9299 3712
rect 9333 3678 9366 3712
rect 26 3644 320 3678
rect 354 3644 379 3678
rect 984 3644 1040 3678
rect 1074 3644 1662 3678
rect 1696 3644 1752 3678
rect 1786 3644 1842 3678
rect 1876 3644 1932 3678
rect 1966 3644 2022 3678
rect 2056 3644 2112 3678
rect 2146 3644 2202 3678
rect 2236 3644 2292 3678
rect 2326 3644 2382 3678
rect 2416 3644 3004 3678
rect 3038 3644 3094 3678
rect 3128 3644 3184 3678
rect 3218 3644 3274 3678
rect 3308 3644 3364 3678
rect 3398 3644 3454 3678
rect 3488 3644 3544 3678
rect 3578 3644 3634 3678
rect 3668 3644 3724 3678
rect 3758 3644 4346 3678
rect 4380 3644 4436 3678
rect 4470 3644 4526 3678
rect 4560 3644 4616 3678
rect 4650 3644 4706 3678
rect 4740 3644 4796 3678
rect 4830 3644 4886 3678
rect 4920 3644 4976 3678
rect 5010 3644 5066 3678
rect 5100 3644 5688 3678
rect 5722 3644 5778 3678
rect 5812 3644 5868 3678
rect 5902 3644 5958 3678
rect 5992 3644 6048 3678
rect 6082 3644 6138 3678
rect 6172 3644 6228 3678
rect 6262 3644 6318 3678
rect 6352 3644 6408 3678
rect 6442 3644 7030 3678
rect 7064 3644 7120 3678
rect 7154 3644 7210 3678
rect 7244 3644 7300 3678
rect 7334 3644 7390 3678
rect 7424 3644 7480 3678
rect 7514 3644 7570 3678
rect 7604 3644 7660 3678
rect 7694 3644 7750 3678
rect 7784 3644 8372 3678
rect 8406 3644 8462 3678
rect 8496 3644 8552 3678
rect 8586 3644 8642 3678
rect 8676 3644 8732 3678
rect 8766 3644 8822 3678
rect 8856 3644 8912 3678
rect 8946 3644 9002 3678
rect 9036 3644 9092 3678
rect 9126 3644 9366 3678
rect 26 3639 379 3644
rect 965 3639 9366 3644
rect 26 3625 9366 3639
rect 26 3622 261 3625
rect 26 3588 60 3622
rect 94 3621 261 3622
rect 94 3588 208 3621
rect 26 3587 208 3588
rect 242 3587 261 3621
rect 26 3532 261 3587
rect 1079 3622 1603 3625
rect 1079 3602 1247 3622
rect 1079 3568 1098 3602
rect 1132 3588 1247 3602
rect 1281 3588 1402 3622
rect 1436 3621 1603 3622
rect 1436 3588 1550 3621
rect 1132 3587 1550 3588
rect 1584 3587 1603 3621
rect 1132 3568 1603 3587
rect 26 3498 60 3532
rect 94 3531 261 3532
rect 94 3498 208 3531
rect 26 3497 208 3498
rect 242 3497 261 3531
rect 26 3442 261 3497
rect 26 3408 60 3442
rect 94 3441 261 3442
rect 94 3408 208 3441
rect 26 3407 208 3408
rect 242 3407 261 3441
rect 26 3352 261 3407
rect 26 3318 60 3352
rect 94 3351 261 3352
rect 94 3318 208 3351
rect 26 3317 208 3318
rect 242 3317 261 3351
rect 26 3262 261 3317
rect 26 3228 60 3262
rect 94 3261 261 3262
rect 94 3228 208 3261
rect 26 3227 208 3228
rect 242 3227 261 3261
rect 26 3172 261 3227
rect 26 3138 60 3172
rect 94 3171 261 3172
rect 94 3138 208 3171
rect 26 3137 208 3138
rect 242 3137 261 3171
rect 26 3082 261 3137
rect 26 3048 60 3082
rect 94 3081 261 3082
rect 94 3048 208 3081
rect 26 3047 208 3048
rect 242 3047 261 3081
rect 26 2992 261 3047
rect 26 2958 60 2992
rect 94 2991 261 2992
rect 94 2958 208 2991
rect 26 2957 208 2958
rect 242 2957 261 2991
rect 26 2902 261 2957
rect 26 2868 60 2902
rect 94 2901 261 2902
rect 94 2868 208 2901
rect 26 2867 208 2868
rect 242 2867 261 2901
rect 323 3504 1017 3563
rect 323 3470 384 3504
rect 418 3470 474 3504
rect 508 3470 564 3504
rect 598 3470 654 3504
rect 688 3470 744 3504
rect 778 3470 834 3504
rect 868 3470 924 3504
rect 958 3470 1017 3504
rect 323 3414 1017 3470
rect 323 3380 384 3414
rect 418 3380 474 3414
rect 508 3380 564 3414
rect 598 3380 654 3414
rect 688 3380 744 3414
rect 778 3380 834 3414
rect 868 3380 924 3414
rect 958 3380 1017 3414
rect 323 3324 1017 3380
rect 323 3290 384 3324
rect 418 3290 474 3324
rect 508 3290 564 3324
rect 598 3290 654 3324
rect 688 3290 744 3324
rect 778 3290 834 3324
rect 868 3290 924 3324
rect 958 3290 1017 3324
rect 323 3234 1017 3290
rect 323 3200 384 3234
rect 418 3200 474 3234
rect 508 3200 564 3234
rect 598 3200 654 3234
rect 688 3200 744 3234
rect 778 3200 834 3234
rect 868 3200 924 3234
rect 958 3200 1017 3234
rect 323 3144 1017 3200
rect 323 3110 384 3144
rect 418 3110 474 3144
rect 508 3110 564 3144
rect 598 3110 654 3144
rect 688 3110 744 3144
rect 778 3110 834 3144
rect 868 3110 924 3144
rect 958 3110 1017 3144
rect 323 3054 1017 3110
rect 323 3020 384 3054
rect 418 3020 474 3054
rect 508 3020 564 3054
rect 598 3020 654 3054
rect 688 3020 744 3054
rect 778 3020 834 3054
rect 868 3020 924 3054
rect 958 3020 1017 3054
rect 323 2964 1017 3020
rect 323 2930 384 2964
rect 418 2930 474 2964
rect 508 2930 564 2964
rect 598 2930 654 2964
rect 688 2930 744 2964
rect 778 2930 834 2964
rect 868 2930 924 2964
rect 958 2930 1017 2964
rect 323 2869 1017 2930
rect 1079 3532 1603 3568
rect 2421 3622 2945 3625
rect 2421 3602 2589 3622
rect 2421 3568 2440 3602
rect 2474 3588 2589 3602
rect 2623 3588 2744 3622
rect 2778 3621 2945 3622
rect 2778 3588 2892 3621
rect 2474 3587 2892 3588
rect 2926 3587 2945 3621
rect 2474 3568 2945 3587
rect 1079 3512 1247 3532
rect 1079 3478 1098 3512
rect 1132 3498 1247 3512
rect 1281 3498 1402 3532
rect 1436 3531 1603 3532
rect 1436 3498 1550 3531
rect 1132 3497 1550 3498
rect 1584 3497 1603 3531
rect 1132 3478 1603 3497
rect 1079 3442 1603 3478
rect 1079 3422 1247 3442
rect 1079 3388 1098 3422
rect 1132 3408 1247 3422
rect 1281 3408 1402 3442
rect 1436 3441 1603 3442
rect 1436 3408 1550 3441
rect 1132 3407 1550 3408
rect 1584 3407 1603 3441
rect 1132 3388 1603 3407
rect 1079 3352 1603 3388
rect 1079 3332 1247 3352
rect 1079 3298 1098 3332
rect 1132 3318 1247 3332
rect 1281 3318 1402 3352
rect 1436 3351 1603 3352
rect 1436 3318 1550 3351
rect 1132 3317 1550 3318
rect 1584 3317 1603 3351
rect 1132 3298 1603 3317
rect 1079 3262 1603 3298
rect 1079 3242 1247 3262
rect 1079 3208 1098 3242
rect 1132 3228 1247 3242
rect 1281 3228 1402 3262
rect 1436 3261 1603 3262
rect 1436 3228 1550 3261
rect 1132 3227 1550 3228
rect 1584 3227 1603 3261
rect 1132 3208 1603 3227
rect 1079 3172 1603 3208
rect 1079 3152 1247 3172
rect 1079 3118 1098 3152
rect 1132 3138 1247 3152
rect 1281 3138 1402 3172
rect 1436 3171 1603 3172
rect 1436 3138 1550 3171
rect 1132 3137 1550 3138
rect 1584 3137 1603 3171
rect 1132 3118 1603 3137
rect 1079 3082 1603 3118
rect 1079 3062 1247 3082
rect 1079 3028 1098 3062
rect 1132 3048 1247 3062
rect 1281 3048 1402 3082
rect 1436 3081 1603 3082
rect 1436 3048 1550 3081
rect 1132 3047 1550 3048
rect 1584 3047 1603 3081
rect 1132 3028 1603 3047
rect 1079 2992 1603 3028
rect 1079 2972 1247 2992
rect 1079 2938 1098 2972
rect 1132 2958 1247 2972
rect 1281 2958 1402 2992
rect 1436 2991 1603 2992
rect 1436 2958 1550 2991
rect 1132 2957 1550 2958
rect 1584 2957 1603 2991
rect 1132 2938 1603 2957
rect 1079 2902 1603 2938
rect 1079 2882 1247 2902
rect 26 2812 261 2867
rect 26 2778 60 2812
rect 94 2807 261 2812
rect 1079 2848 1098 2882
rect 1132 2868 1247 2882
rect 1281 2868 1402 2902
rect 1436 2901 1603 2902
rect 1436 2868 1550 2901
rect 1132 2867 1550 2868
rect 1584 2867 1603 2901
rect 1665 3504 2359 3563
rect 1665 3470 1726 3504
rect 1760 3470 1816 3504
rect 1850 3470 1906 3504
rect 1940 3470 1996 3504
rect 2030 3470 2086 3504
rect 2120 3470 2176 3504
rect 2210 3470 2266 3504
rect 2300 3470 2359 3504
rect 1665 3414 2359 3470
rect 1665 3380 1726 3414
rect 1760 3380 1816 3414
rect 1850 3380 1906 3414
rect 1940 3380 1996 3414
rect 2030 3380 2086 3414
rect 2120 3380 2176 3414
rect 2210 3380 2266 3414
rect 2300 3380 2359 3414
rect 1665 3324 2359 3380
rect 1665 3290 1726 3324
rect 1760 3290 1816 3324
rect 1850 3290 1906 3324
rect 1940 3290 1996 3324
rect 2030 3290 2086 3324
rect 2120 3290 2176 3324
rect 2210 3290 2266 3324
rect 2300 3290 2359 3324
rect 1665 3234 2359 3290
rect 1665 3200 1726 3234
rect 1760 3200 1816 3234
rect 1850 3200 1906 3234
rect 1940 3200 1996 3234
rect 2030 3200 2086 3234
rect 2120 3200 2176 3234
rect 2210 3200 2266 3234
rect 2300 3200 2359 3234
rect 1665 3144 2359 3200
rect 1665 3110 1726 3144
rect 1760 3110 1816 3144
rect 1850 3110 1906 3144
rect 1940 3110 1996 3144
rect 2030 3110 2086 3144
rect 2120 3110 2176 3144
rect 2210 3110 2266 3144
rect 2300 3110 2359 3144
rect 1665 3054 2359 3110
rect 1665 3020 1726 3054
rect 1760 3020 1816 3054
rect 1850 3020 1906 3054
rect 1940 3020 1996 3054
rect 2030 3020 2086 3054
rect 2120 3020 2176 3054
rect 2210 3020 2266 3054
rect 2300 3020 2359 3054
rect 1665 2964 2359 3020
rect 1665 2930 1726 2964
rect 1760 2930 1816 2964
rect 1850 2930 1906 2964
rect 1940 2930 1996 2964
rect 2030 2930 2086 2964
rect 2120 2930 2176 2964
rect 2210 2930 2266 2964
rect 2300 2930 2359 2964
rect 1665 2869 2359 2930
rect 2421 3532 2945 3568
rect 3763 3622 4287 3625
rect 3763 3602 3931 3622
rect 3763 3568 3782 3602
rect 3816 3588 3931 3602
rect 3965 3588 4086 3622
rect 4120 3621 4287 3622
rect 4120 3588 4234 3621
rect 3816 3587 4234 3588
rect 4268 3587 4287 3621
rect 3816 3568 4287 3587
rect 2421 3512 2589 3532
rect 2421 3478 2440 3512
rect 2474 3498 2589 3512
rect 2623 3498 2744 3532
rect 2778 3531 2945 3532
rect 2778 3498 2892 3531
rect 2474 3497 2892 3498
rect 2926 3497 2945 3531
rect 2474 3478 2945 3497
rect 2421 3442 2945 3478
rect 2421 3422 2589 3442
rect 2421 3388 2440 3422
rect 2474 3408 2589 3422
rect 2623 3408 2744 3442
rect 2778 3441 2945 3442
rect 2778 3408 2892 3441
rect 2474 3407 2892 3408
rect 2926 3407 2945 3441
rect 2474 3388 2945 3407
rect 2421 3352 2945 3388
rect 2421 3332 2589 3352
rect 2421 3298 2440 3332
rect 2474 3318 2589 3332
rect 2623 3318 2744 3352
rect 2778 3351 2945 3352
rect 2778 3318 2892 3351
rect 2474 3317 2892 3318
rect 2926 3317 2945 3351
rect 2474 3298 2945 3317
rect 2421 3262 2945 3298
rect 2421 3242 2589 3262
rect 2421 3208 2440 3242
rect 2474 3228 2589 3242
rect 2623 3228 2744 3262
rect 2778 3261 2945 3262
rect 2778 3228 2892 3261
rect 2474 3227 2892 3228
rect 2926 3227 2945 3261
rect 2474 3208 2945 3227
rect 2421 3172 2945 3208
rect 2421 3152 2589 3172
rect 2421 3118 2440 3152
rect 2474 3138 2589 3152
rect 2623 3138 2744 3172
rect 2778 3171 2945 3172
rect 2778 3138 2892 3171
rect 2474 3137 2892 3138
rect 2926 3137 2945 3171
rect 2474 3118 2945 3137
rect 2421 3082 2945 3118
rect 2421 3062 2589 3082
rect 2421 3028 2440 3062
rect 2474 3048 2589 3062
rect 2623 3048 2744 3082
rect 2778 3081 2945 3082
rect 2778 3048 2892 3081
rect 2474 3047 2892 3048
rect 2926 3047 2945 3081
rect 2474 3028 2945 3047
rect 2421 2992 2945 3028
rect 2421 2972 2589 2992
rect 2421 2938 2440 2972
rect 2474 2958 2589 2972
rect 2623 2958 2744 2992
rect 2778 2991 2945 2992
rect 2778 2958 2892 2991
rect 2474 2957 2892 2958
rect 2926 2957 2945 2991
rect 2474 2938 2945 2957
rect 2421 2902 2945 2938
rect 2421 2882 2589 2902
rect 1132 2848 1603 2867
rect 1079 2812 1603 2848
rect 1079 2807 1247 2812
rect 94 2788 1247 2807
rect 94 2778 286 2788
rect 26 2754 286 2778
rect 320 2754 376 2788
rect 410 2754 466 2788
rect 500 2754 556 2788
rect 590 2754 646 2788
rect 680 2754 736 2788
rect 770 2754 826 2788
rect 860 2754 916 2788
rect 950 2754 1006 2788
rect 1040 2778 1247 2788
rect 1281 2778 1402 2812
rect 1436 2807 1603 2812
rect 2421 2848 2440 2882
rect 2474 2868 2589 2882
rect 2623 2868 2744 2902
rect 2778 2901 2945 2902
rect 2778 2868 2892 2901
rect 2474 2867 2892 2868
rect 2926 2867 2945 2901
rect 3007 3504 3701 3563
rect 3007 3470 3068 3504
rect 3102 3470 3158 3504
rect 3192 3470 3248 3504
rect 3282 3470 3338 3504
rect 3372 3470 3428 3504
rect 3462 3470 3518 3504
rect 3552 3470 3608 3504
rect 3642 3470 3701 3504
rect 3007 3414 3701 3470
rect 3007 3380 3068 3414
rect 3102 3380 3158 3414
rect 3192 3380 3248 3414
rect 3282 3380 3338 3414
rect 3372 3380 3428 3414
rect 3462 3380 3518 3414
rect 3552 3380 3608 3414
rect 3642 3380 3701 3414
rect 3007 3324 3701 3380
rect 3007 3290 3068 3324
rect 3102 3290 3158 3324
rect 3192 3290 3248 3324
rect 3282 3290 3338 3324
rect 3372 3290 3428 3324
rect 3462 3290 3518 3324
rect 3552 3290 3608 3324
rect 3642 3290 3701 3324
rect 3007 3234 3701 3290
rect 3007 3200 3068 3234
rect 3102 3200 3158 3234
rect 3192 3200 3248 3234
rect 3282 3200 3338 3234
rect 3372 3200 3428 3234
rect 3462 3200 3518 3234
rect 3552 3200 3608 3234
rect 3642 3200 3701 3234
rect 3007 3144 3701 3200
rect 3007 3110 3068 3144
rect 3102 3110 3158 3144
rect 3192 3110 3248 3144
rect 3282 3110 3338 3144
rect 3372 3110 3428 3144
rect 3462 3110 3518 3144
rect 3552 3110 3608 3144
rect 3642 3110 3701 3144
rect 3007 3054 3701 3110
rect 3007 3020 3068 3054
rect 3102 3020 3158 3054
rect 3192 3020 3248 3054
rect 3282 3020 3338 3054
rect 3372 3020 3428 3054
rect 3462 3020 3518 3054
rect 3552 3020 3608 3054
rect 3642 3020 3701 3054
rect 3007 2964 3701 3020
rect 3007 2930 3068 2964
rect 3102 2930 3158 2964
rect 3192 2930 3248 2964
rect 3282 2930 3338 2964
rect 3372 2930 3428 2964
rect 3462 2930 3518 2964
rect 3552 2930 3608 2964
rect 3642 2930 3701 2964
rect 3007 2869 3701 2930
rect 3763 3532 4287 3568
rect 5105 3622 5629 3625
rect 5105 3602 5273 3622
rect 5105 3568 5124 3602
rect 5158 3588 5273 3602
rect 5307 3588 5428 3622
rect 5462 3621 5629 3622
rect 5462 3588 5576 3621
rect 5158 3587 5576 3588
rect 5610 3587 5629 3621
rect 5158 3568 5629 3587
rect 3763 3512 3931 3532
rect 3763 3478 3782 3512
rect 3816 3498 3931 3512
rect 3965 3498 4086 3532
rect 4120 3531 4287 3532
rect 4120 3498 4234 3531
rect 3816 3497 4234 3498
rect 4268 3497 4287 3531
rect 3816 3478 4287 3497
rect 3763 3442 4287 3478
rect 3763 3422 3931 3442
rect 3763 3388 3782 3422
rect 3816 3408 3931 3422
rect 3965 3408 4086 3442
rect 4120 3441 4287 3442
rect 4120 3408 4234 3441
rect 3816 3407 4234 3408
rect 4268 3407 4287 3441
rect 3816 3388 4287 3407
rect 3763 3352 4287 3388
rect 3763 3332 3931 3352
rect 3763 3298 3782 3332
rect 3816 3318 3931 3332
rect 3965 3318 4086 3352
rect 4120 3351 4287 3352
rect 4120 3318 4234 3351
rect 3816 3317 4234 3318
rect 4268 3317 4287 3351
rect 3816 3298 4287 3317
rect 3763 3262 4287 3298
rect 3763 3242 3931 3262
rect 3763 3208 3782 3242
rect 3816 3228 3931 3242
rect 3965 3228 4086 3262
rect 4120 3261 4287 3262
rect 4120 3228 4234 3261
rect 3816 3227 4234 3228
rect 4268 3227 4287 3261
rect 3816 3208 4287 3227
rect 3763 3172 4287 3208
rect 3763 3152 3931 3172
rect 3763 3118 3782 3152
rect 3816 3138 3931 3152
rect 3965 3138 4086 3172
rect 4120 3171 4287 3172
rect 4120 3138 4234 3171
rect 3816 3137 4234 3138
rect 4268 3137 4287 3171
rect 3816 3118 4287 3137
rect 3763 3082 4287 3118
rect 3763 3062 3931 3082
rect 3763 3028 3782 3062
rect 3816 3048 3931 3062
rect 3965 3048 4086 3082
rect 4120 3081 4287 3082
rect 4120 3048 4234 3081
rect 3816 3047 4234 3048
rect 4268 3047 4287 3081
rect 3816 3028 4287 3047
rect 3763 2992 4287 3028
rect 3763 2972 3931 2992
rect 3763 2938 3782 2972
rect 3816 2958 3931 2972
rect 3965 2958 4086 2992
rect 4120 2991 4287 2992
rect 4120 2958 4234 2991
rect 3816 2957 4234 2958
rect 4268 2957 4287 2991
rect 3816 2938 4287 2957
rect 3763 2902 4287 2938
rect 3763 2882 3931 2902
rect 2474 2848 2945 2867
rect 2421 2812 2945 2848
rect 2421 2807 2589 2812
rect 1436 2788 2589 2807
rect 1436 2778 1628 2788
rect 1040 2754 1628 2778
rect 1662 2754 1718 2788
rect 1752 2754 1808 2788
rect 1842 2754 1898 2788
rect 1932 2754 1988 2788
rect 2022 2754 2078 2788
rect 2112 2754 2168 2788
rect 2202 2754 2258 2788
rect 2292 2754 2348 2788
rect 2382 2778 2589 2788
rect 2623 2778 2744 2812
rect 2778 2807 2945 2812
rect 3763 2848 3782 2882
rect 3816 2868 3931 2882
rect 3965 2868 4086 2902
rect 4120 2901 4287 2902
rect 4120 2868 4234 2901
rect 3816 2867 4234 2868
rect 4268 2867 4287 2901
rect 4349 3504 5043 3563
rect 4349 3470 4410 3504
rect 4444 3470 4500 3504
rect 4534 3470 4590 3504
rect 4624 3470 4680 3504
rect 4714 3470 4770 3504
rect 4804 3470 4860 3504
rect 4894 3470 4950 3504
rect 4984 3470 5043 3504
rect 4349 3414 5043 3470
rect 4349 3380 4410 3414
rect 4444 3380 4500 3414
rect 4534 3380 4590 3414
rect 4624 3380 4680 3414
rect 4714 3380 4770 3414
rect 4804 3380 4860 3414
rect 4894 3380 4950 3414
rect 4984 3380 5043 3414
rect 4349 3324 5043 3380
rect 4349 3290 4410 3324
rect 4444 3290 4500 3324
rect 4534 3290 4590 3324
rect 4624 3290 4680 3324
rect 4714 3290 4770 3324
rect 4804 3290 4860 3324
rect 4894 3290 4950 3324
rect 4984 3290 5043 3324
rect 4349 3234 5043 3290
rect 4349 3200 4410 3234
rect 4444 3200 4500 3234
rect 4534 3200 4590 3234
rect 4624 3200 4680 3234
rect 4714 3200 4770 3234
rect 4804 3200 4860 3234
rect 4894 3200 4950 3234
rect 4984 3200 5043 3234
rect 4349 3144 5043 3200
rect 4349 3110 4410 3144
rect 4444 3110 4500 3144
rect 4534 3110 4590 3144
rect 4624 3110 4680 3144
rect 4714 3110 4770 3144
rect 4804 3110 4860 3144
rect 4894 3110 4950 3144
rect 4984 3110 5043 3144
rect 4349 3054 5043 3110
rect 4349 3020 4410 3054
rect 4444 3020 4500 3054
rect 4534 3020 4590 3054
rect 4624 3020 4680 3054
rect 4714 3020 4770 3054
rect 4804 3020 4860 3054
rect 4894 3020 4950 3054
rect 4984 3020 5043 3054
rect 4349 2964 5043 3020
rect 4349 2930 4410 2964
rect 4444 2930 4500 2964
rect 4534 2930 4590 2964
rect 4624 2930 4680 2964
rect 4714 2930 4770 2964
rect 4804 2930 4860 2964
rect 4894 2930 4950 2964
rect 4984 2930 5043 2964
rect 4349 2869 5043 2930
rect 5105 3532 5629 3568
rect 6447 3622 6971 3625
rect 6447 3602 6615 3622
rect 6447 3568 6466 3602
rect 6500 3588 6615 3602
rect 6649 3588 6770 3622
rect 6804 3621 6971 3622
rect 6804 3588 6918 3621
rect 6500 3587 6918 3588
rect 6952 3587 6971 3621
rect 6500 3568 6971 3587
rect 5105 3512 5273 3532
rect 5105 3478 5124 3512
rect 5158 3498 5273 3512
rect 5307 3498 5428 3532
rect 5462 3531 5629 3532
rect 5462 3498 5576 3531
rect 5158 3497 5576 3498
rect 5610 3497 5629 3531
rect 5158 3478 5629 3497
rect 5105 3442 5629 3478
rect 5105 3422 5273 3442
rect 5105 3388 5124 3422
rect 5158 3408 5273 3422
rect 5307 3408 5428 3442
rect 5462 3441 5629 3442
rect 5462 3408 5576 3441
rect 5158 3407 5576 3408
rect 5610 3407 5629 3441
rect 5158 3388 5629 3407
rect 5105 3352 5629 3388
rect 5105 3332 5273 3352
rect 5105 3298 5124 3332
rect 5158 3318 5273 3332
rect 5307 3318 5428 3352
rect 5462 3351 5629 3352
rect 5462 3318 5576 3351
rect 5158 3317 5576 3318
rect 5610 3317 5629 3351
rect 5158 3298 5629 3317
rect 5105 3262 5629 3298
rect 5105 3242 5273 3262
rect 5105 3208 5124 3242
rect 5158 3228 5273 3242
rect 5307 3228 5428 3262
rect 5462 3261 5629 3262
rect 5462 3228 5576 3261
rect 5158 3227 5576 3228
rect 5610 3227 5629 3261
rect 5158 3208 5629 3227
rect 5105 3172 5629 3208
rect 5105 3152 5273 3172
rect 5105 3118 5124 3152
rect 5158 3138 5273 3152
rect 5307 3138 5428 3172
rect 5462 3171 5629 3172
rect 5462 3138 5576 3171
rect 5158 3137 5576 3138
rect 5610 3137 5629 3171
rect 5158 3118 5629 3137
rect 5105 3082 5629 3118
rect 5105 3062 5273 3082
rect 5105 3028 5124 3062
rect 5158 3048 5273 3062
rect 5307 3048 5428 3082
rect 5462 3081 5629 3082
rect 5462 3048 5576 3081
rect 5158 3047 5576 3048
rect 5610 3047 5629 3081
rect 5158 3028 5629 3047
rect 5105 2992 5629 3028
rect 5105 2972 5273 2992
rect 5105 2938 5124 2972
rect 5158 2958 5273 2972
rect 5307 2958 5428 2992
rect 5462 2991 5629 2992
rect 5462 2958 5576 2991
rect 5158 2957 5576 2958
rect 5610 2957 5629 2991
rect 5158 2938 5629 2957
rect 5105 2902 5629 2938
rect 5105 2882 5273 2902
rect 3816 2848 4287 2867
rect 3763 2812 4287 2848
rect 3763 2807 3931 2812
rect 2778 2788 3931 2807
rect 2778 2778 2970 2788
rect 2382 2754 2970 2778
rect 3004 2754 3060 2788
rect 3094 2754 3150 2788
rect 3184 2754 3240 2788
rect 3274 2754 3330 2788
rect 3364 2754 3420 2788
rect 3454 2754 3510 2788
rect 3544 2754 3600 2788
rect 3634 2754 3690 2788
rect 3724 2778 3931 2788
rect 3965 2778 4086 2812
rect 4120 2807 4287 2812
rect 5105 2848 5124 2882
rect 5158 2868 5273 2882
rect 5307 2868 5428 2902
rect 5462 2901 5629 2902
rect 5462 2868 5576 2901
rect 5158 2867 5576 2868
rect 5610 2867 5629 2901
rect 5691 3504 6385 3563
rect 5691 3470 5752 3504
rect 5786 3470 5842 3504
rect 5876 3470 5932 3504
rect 5966 3470 6022 3504
rect 6056 3470 6112 3504
rect 6146 3470 6202 3504
rect 6236 3470 6292 3504
rect 6326 3470 6385 3504
rect 5691 3414 6385 3470
rect 5691 3380 5752 3414
rect 5786 3380 5842 3414
rect 5876 3380 5932 3414
rect 5966 3380 6022 3414
rect 6056 3380 6112 3414
rect 6146 3380 6202 3414
rect 6236 3380 6292 3414
rect 6326 3380 6385 3414
rect 5691 3324 6385 3380
rect 5691 3290 5752 3324
rect 5786 3290 5842 3324
rect 5876 3290 5932 3324
rect 5966 3290 6022 3324
rect 6056 3290 6112 3324
rect 6146 3290 6202 3324
rect 6236 3290 6292 3324
rect 6326 3290 6385 3324
rect 5691 3234 6385 3290
rect 5691 3200 5752 3234
rect 5786 3200 5842 3234
rect 5876 3200 5932 3234
rect 5966 3200 6022 3234
rect 6056 3200 6112 3234
rect 6146 3200 6202 3234
rect 6236 3200 6292 3234
rect 6326 3200 6385 3234
rect 5691 3144 6385 3200
rect 5691 3110 5752 3144
rect 5786 3110 5842 3144
rect 5876 3110 5932 3144
rect 5966 3110 6022 3144
rect 6056 3110 6112 3144
rect 6146 3110 6202 3144
rect 6236 3110 6292 3144
rect 6326 3110 6385 3144
rect 5691 3054 6385 3110
rect 5691 3020 5752 3054
rect 5786 3020 5842 3054
rect 5876 3020 5932 3054
rect 5966 3020 6022 3054
rect 6056 3020 6112 3054
rect 6146 3020 6202 3054
rect 6236 3020 6292 3054
rect 6326 3020 6385 3054
rect 5691 2964 6385 3020
rect 5691 2930 5752 2964
rect 5786 2930 5842 2964
rect 5876 2930 5932 2964
rect 5966 2930 6022 2964
rect 6056 2930 6112 2964
rect 6146 2930 6202 2964
rect 6236 2930 6292 2964
rect 6326 2930 6385 2964
rect 5691 2869 6385 2930
rect 6447 3532 6971 3568
rect 7789 3622 8313 3625
rect 7789 3602 7957 3622
rect 7789 3568 7808 3602
rect 7842 3588 7957 3602
rect 7991 3588 8112 3622
rect 8146 3621 8313 3622
rect 8146 3588 8260 3621
rect 7842 3587 8260 3588
rect 8294 3587 8313 3621
rect 7842 3568 8313 3587
rect 6447 3512 6615 3532
rect 6447 3478 6466 3512
rect 6500 3498 6615 3512
rect 6649 3498 6770 3532
rect 6804 3531 6971 3532
rect 6804 3498 6918 3531
rect 6500 3497 6918 3498
rect 6952 3497 6971 3531
rect 6500 3478 6971 3497
rect 6447 3442 6971 3478
rect 6447 3422 6615 3442
rect 6447 3388 6466 3422
rect 6500 3408 6615 3422
rect 6649 3408 6770 3442
rect 6804 3441 6971 3442
rect 6804 3408 6918 3441
rect 6500 3407 6918 3408
rect 6952 3407 6971 3441
rect 6500 3388 6971 3407
rect 6447 3352 6971 3388
rect 6447 3332 6615 3352
rect 6447 3298 6466 3332
rect 6500 3318 6615 3332
rect 6649 3318 6770 3352
rect 6804 3351 6971 3352
rect 6804 3318 6918 3351
rect 6500 3317 6918 3318
rect 6952 3317 6971 3351
rect 6500 3298 6971 3317
rect 6447 3262 6971 3298
rect 6447 3242 6615 3262
rect 6447 3208 6466 3242
rect 6500 3228 6615 3242
rect 6649 3228 6770 3262
rect 6804 3261 6971 3262
rect 6804 3228 6918 3261
rect 6500 3227 6918 3228
rect 6952 3227 6971 3261
rect 6500 3208 6971 3227
rect 6447 3172 6971 3208
rect 6447 3152 6615 3172
rect 6447 3118 6466 3152
rect 6500 3138 6615 3152
rect 6649 3138 6770 3172
rect 6804 3171 6971 3172
rect 6804 3138 6918 3171
rect 6500 3137 6918 3138
rect 6952 3137 6971 3171
rect 6500 3118 6971 3137
rect 6447 3082 6971 3118
rect 6447 3062 6615 3082
rect 6447 3028 6466 3062
rect 6500 3048 6615 3062
rect 6649 3048 6770 3082
rect 6804 3081 6971 3082
rect 6804 3048 6918 3081
rect 6500 3047 6918 3048
rect 6952 3047 6971 3081
rect 6500 3028 6971 3047
rect 6447 2992 6971 3028
rect 6447 2972 6615 2992
rect 6447 2938 6466 2972
rect 6500 2958 6615 2972
rect 6649 2958 6770 2992
rect 6804 2991 6971 2992
rect 6804 2958 6918 2991
rect 6500 2957 6918 2958
rect 6952 2957 6971 2991
rect 6500 2938 6971 2957
rect 6447 2902 6971 2938
rect 6447 2882 6615 2902
rect 5158 2848 5629 2867
rect 5105 2812 5629 2848
rect 5105 2807 5273 2812
rect 4120 2788 5273 2807
rect 4120 2778 4312 2788
rect 3724 2754 4312 2778
rect 4346 2754 4402 2788
rect 4436 2754 4492 2788
rect 4526 2754 4582 2788
rect 4616 2754 4672 2788
rect 4706 2754 4762 2788
rect 4796 2754 4852 2788
rect 4886 2754 4942 2788
rect 4976 2754 5032 2788
rect 5066 2778 5273 2788
rect 5307 2778 5428 2812
rect 5462 2807 5629 2812
rect 6447 2848 6466 2882
rect 6500 2868 6615 2882
rect 6649 2868 6770 2902
rect 6804 2901 6971 2902
rect 6804 2868 6918 2901
rect 6500 2867 6918 2868
rect 6952 2867 6971 2901
rect 7033 3504 7727 3563
rect 7033 3470 7094 3504
rect 7128 3470 7184 3504
rect 7218 3470 7274 3504
rect 7308 3470 7364 3504
rect 7398 3470 7454 3504
rect 7488 3470 7544 3504
rect 7578 3470 7634 3504
rect 7668 3470 7727 3504
rect 7033 3414 7727 3470
rect 7033 3380 7094 3414
rect 7128 3380 7184 3414
rect 7218 3380 7274 3414
rect 7308 3380 7364 3414
rect 7398 3380 7454 3414
rect 7488 3380 7544 3414
rect 7578 3380 7634 3414
rect 7668 3380 7727 3414
rect 7033 3324 7727 3380
rect 7033 3290 7094 3324
rect 7128 3290 7184 3324
rect 7218 3290 7274 3324
rect 7308 3290 7364 3324
rect 7398 3290 7454 3324
rect 7488 3290 7544 3324
rect 7578 3290 7634 3324
rect 7668 3290 7727 3324
rect 7033 3234 7727 3290
rect 7033 3200 7094 3234
rect 7128 3200 7184 3234
rect 7218 3200 7274 3234
rect 7308 3200 7364 3234
rect 7398 3200 7454 3234
rect 7488 3200 7544 3234
rect 7578 3200 7634 3234
rect 7668 3200 7727 3234
rect 7033 3144 7727 3200
rect 7033 3110 7094 3144
rect 7128 3110 7184 3144
rect 7218 3110 7274 3144
rect 7308 3110 7364 3144
rect 7398 3110 7454 3144
rect 7488 3110 7544 3144
rect 7578 3110 7634 3144
rect 7668 3110 7727 3144
rect 7033 3054 7727 3110
rect 7033 3020 7094 3054
rect 7128 3020 7184 3054
rect 7218 3020 7274 3054
rect 7308 3020 7364 3054
rect 7398 3020 7454 3054
rect 7488 3020 7544 3054
rect 7578 3020 7634 3054
rect 7668 3020 7727 3054
rect 7033 2964 7727 3020
rect 7033 2930 7094 2964
rect 7128 2930 7184 2964
rect 7218 2930 7274 2964
rect 7308 2930 7364 2964
rect 7398 2930 7454 2964
rect 7488 2930 7544 2964
rect 7578 2930 7634 2964
rect 7668 2930 7727 2964
rect 7033 2869 7727 2930
rect 7789 3532 8313 3568
rect 9131 3622 9366 3625
rect 9131 3602 9299 3622
rect 9131 3568 9150 3602
rect 9184 3588 9299 3602
rect 9333 3588 9366 3622
rect 9184 3568 9366 3588
rect 7789 3512 7957 3532
rect 7789 3478 7808 3512
rect 7842 3498 7957 3512
rect 7991 3498 8112 3532
rect 8146 3531 8313 3532
rect 8146 3498 8260 3531
rect 7842 3497 8260 3498
rect 8294 3497 8313 3531
rect 7842 3478 8313 3497
rect 7789 3442 8313 3478
rect 7789 3422 7957 3442
rect 7789 3388 7808 3422
rect 7842 3408 7957 3422
rect 7991 3408 8112 3442
rect 8146 3441 8313 3442
rect 8146 3408 8260 3441
rect 7842 3407 8260 3408
rect 8294 3407 8313 3441
rect 7842 3388 8313 3407
rect 7789 3352 8313 3388
rect 7789 3332 7957 3352
rect 7789 3298 7808 3332
rect 7842 3318 7957 3332
rect 7991 3318 8112 3352
rect 8146 3351 8313 3352
rect 8146 3318 8260 3351
rect 7842 3317 8260 3318
rect 8294 3317 8313 3351
rect 7842 3298 8313 3317
rect 7789 3262 8313 3298
rect 7789 3242 7957 3262
rect 7789 3208 7808 3242
rect 7842 3228 7957 3242
rect 7991 3228 8112 3262
rect 8146 3261 8313 3262
rect 8146 3228 8260 3261
rect 7842 3227 8260 3228
rect 8294 3227 8313 3261
rect 7842 3208 8313 3227
rect 7789 3172 8313 3208
rect 7789 3152 7957 3172
rect 7789 3118 7808 3152
rect 7842 3138 7957 3152
rect 7991 3138 8112 3172
rect 8146 3171 8313 3172
rect 8146 3138 8260 3171
rect 7842 3137 8260 3138
rect 8294 3137 8313 3171
rect 7842 3118 8313 3137
rect 7789 3082 8313 3118
rect 7789 3062 7957 3082
rect 7789 3028 7808 3062
rect 7842 3048 7957 3062
rect 7991 3048 8112 3082
rect 8146 3081 8313 3082
rect 8146 3048 8260 3081
rect 7842 3047 8260 3048
rect 8294 3047 8313 3081
rect 7842 3028 8313 3047
rect 7789 2992 8313 3028
rect 7789 2972 7957 2992
rect 7789 2938 7808 2972
rect 7842 2958 7957 2972
rect 7991 2958 8112 2992
rect 8146 2991 8313 2992
rect 8146 2958 8260 2991
rect 7842 2957 8260 2958
rect 8294 2957 8313 2991
rect 7842 2938 8313 2957
rect 7789 2902 8313 2938
rect 7789 2882 7957 2902
rect 6500 2848 6971 2867
rect 6447 2812 6971 2848
rect 6447 2807 6615 2812
rect 5462 2788 6615 2807
rect 5462 2778 5654 2788
rect 5066 2754 5654 2778
rect 5688 2754 5744 2788
rect 5778 2754 5834 2788
rect 5868 2754 5924 2788
rect 5958 2754 6014 2788
rect 6048 2754 6104 2788
rect 6138 2754 6194 2788
rect 6228 2754 6284 2788
rect 6318 2754 6374 2788
rect 6408 2778 6615 2788
rect 6649 2778 6770 2812
rect 6804 2807 6971 2812
rect 7789 2848 7808 2882
rect 7842 2868 7957 2882
rect 7991 2868 8112 2902
rect 8146 2901 8313 2902
rect 8146 2868 8260 2901
rect 7842 2867 8260 2868
rect 8294 2867 8313 2901
rect 8375 3504 9069 3563
rect 8375 3470 8436 3504
rect 8470 3470 8526 3504
rect 8560 3470 8616 3504
rect 8650 3470 8706 3504
rect 8740 3470 8796 3504
rect 8830 3470 8886 3504
rect 8920 3470 8976 3504
rect 9010 3470 9069 3504
rect 8375 3414 9069 3470
rect 8375 3380 8436 3414
rect 8470 3380 8526 3414
rect 8560 3380 8616 3414
rect 8650 3380 8706 3414
rect 8740 3380 8796 3414
rect 8830 3380 8886 3414
rect 8920 3380 8976 3414
rect 9010 3380 9069 3414
rect 8375 3324 9069 3380
rect 8375 3290 8436 3324
rect 8470 3290 8526 3324
rect 8560 3290 8616 3324
rect 8650 3290 8706 3324
rect 8740 3290 8796 3324
rect 8830 3290 8886 3324
rect 8920 3290 8976 3324
rect 9010 3290 9069 3324
rect 8375 3234 9069 3290
rect 8375 3200 8436 3234
rect 8470 3200 8526 3234
rect 8560 3200 8616 3234
rect 8650 3200 8706 3234
rect 8740 3200 8796 3234
rect 8830 3200 8886 3234
rect 8920 3200 8976 3234
rect 9010 3200 9069 3234
rect 8375 3144 9069 3200
rect 8375 3110 8436 3144
rect 8470 3110 8526 3144
rect 8560 3110 8616 3144
rect 8650 3110 8706 3144
rect 8740 3110 8796 3144
rect 8830 3110 8886 3144
rect 8920 3110 8976 3144
rect 9010 3110 9069 3144
rect 8375 3054 9069 3110
rect 8375 3020 8436 3054
rect 8470 3020 8526 3054
rect 8560 3020 8616 3054
rect 8650 3020 8706 3054
rect 8740 3020 8796 3054
rect 8830 3020 8886 3054
rect 8920 3020 8976 3054
rect 9010 3020 9069 3054
rect 8375 2964 9069 3020
rect 8375 2930 8436 2964
rect 8470 2930 8526 2964
rect 8560 2930 8616 2964
rect 8650 2930 8706 2964
rect 8740 2930 8796 2964
rect 8830 2930 8886 2964
rect 8920 2930 8976 2964
rect 9010 2930 9069 2964
rect 8375 2869 9069 2930
rect 9131 3532 9366 3568
rect 9131 3512 9299 3532
rect 9131 3478 9150 3512
rect 9184 3498 9299 3512
rect 9333 3498 9366 3532
rect 9184 3478 9366 3498
rect 9131 3442 9366 3478
rect 9131 3422 9299 3442
rect 9131 3388 9150 3422
rect 9184 3408 9299 3422
rect 9333 3408 9366 3442
rect 9184 3388 9366 3408
rect 9131 3352 9366 3388
rect 9131 3332 9299 3352
rect 9131 3298 9150 3332
rect 9184 3318 9299 3332
rect 9333 3318 9366 3352
rect 9184 3298 9366 3318
rect 9131 3262 9366 3298
rect 9131 3242 9299 3262
rect 9131 3208 9150 3242
rect 9184 3228 9299 3242
rect 9333 3228 9366 3262
rect 9184 3208 9366 3228
rect 9131 3172 9366 3208
rect 9131 3152 9299 3172
rect 9131 3118 9150 3152
rect 9184 3138 9299 3152
rect 9333 3138 9366 3172
rect 9184 3118 9366 3138
rect 9131 3082 9366 3118
rect 9131 3062 9299 3082
rect 9131 3028 9150 3062
rect 9184 3048 9299 3062
rect 9333 3048 9366 3082
rect 9184 3028 9366 3048
rect 9131 2992 9366 3028
rect 9131 2972 9299 2992
rect 9131 2938 9150 2972
rect 9184 2958 9299 2972
rect 9333 2958 9366 2992
rect 9184 2938 9366 2958
rect 9131 2902 9366 2938
rect 9131 2882 9299 2902
rect 7842 2848 8313 2867
rect 7789 2812 8313 2848
rect 7789 2807 7957 2812
rect 6804 2788 7957 2807
rect 6804 2778 6996 2788
rect 6408 2754 6996 2778
rect 7030 2754 7086 2788
rect 7120 2754 7176 2788
rect 7210 2754 7266 2788
rect 7300 2754 7356 2788
rect 7390 2754 7446 2788
rect 7480 2754 7536 2788
rect 7570 2754 7626 2788
rect 7660 2754 7716 2788
rect 7750 2778 7957 2788
rect 7991 2778 8112 2812
rect 8146 2807 8313 2812
rect 9131 2848 9150 2882
rect 9184 2868 9299 2882
rect 9333 2868 9366 2902
rect 9184 2848 9366 2868
rect 9131 2812 9366 2848
rect 9131 2807 9299 2812
rect 8146 2788 9299 2807
rect 8146 2778 8338 2788
rect 7750 2754 8338 2778
rect 8372 2754 8428 2788
rect 8462 2754 8518 2788
rect 8552 2754 8608 2788
rect 8642 2754 8698 2788
rect 8732 2754 8788 2788
rect 8822 2754 8878 2788
rect 8912 2754 8968 2788
rect 9002 2754 9058 2788
rect 9092 2778 9299 2788
rect 9333 2778 9366 2812
rect 9092 2754 9366 2778
rect 26 2722 9366 2754
rect 26 2688 60 2722
rect 94 2688 1247 2722
rect 1281 2688 1402 2722
rect 1436 2688 2589 2722
rect 2623 2688 2744 2722
rect 2778 2688 3931 2722
rect 3965 2688 4086 2722
rect 4120 2688 5273 2722
rect 5307 2688 5428 2722
rect 5462 2688 6615 2722
rect 6649 2688 6770 2722
rect 6804 2688 7957 2722
rect 7991 2688 8112 2722
rect 8146 2688 9299 2722
rect 9333 2688 9366 2722
rect 26 2638 9366 2688
rect 26 2604 156 2638
rect 190 2604 246 2638
rect 280 2604 336 2638
rect 370 2604 426 2638
rect 460 2604 516 2638
rect 550 2604 606 2638
rect 640 2604 696 2638
rect 730 2604 786 2638
rect 820 2604 876 2638
rect 910 2604 966 2638
rect 1000 2604 1056 2638
rect 1090 2604 1146 2638
rect 1180 2604 1498 2638
rect 1532 2604 1588 2638
rect 1622 2604 1678 2638
rect 1712 2604 1768 2638
rect 1802 2604 1858 2638
rect 1892 2604 1948 2638
rect 1982 2604 2038 2638
rect 2072 2604 2128 2638
rect 2162 2604 2218 2638
rect 2252 2604 2308 2638
rect 2342 2604 2398 2638
rect 2432 2604 2488 2638
rect 2522 2604 2840 2638
rect 2874 2604 2930 2638
rect 2964 2604 3020 2638
rect 3054 2604 3110 2638
rect 3144 2604 3200 2638
rect 3234 2604 3290 2638
rect 3324 2604 3380 2638
rect 3414 2604 3470 2638
rect 3504 2604 3560 2638
rect 3594 2604 3650 2638
rect 3684 2604 3740 2638
rect 3774 2604 3830 2638
rect 3864 2604 4182 2638
rect 4216 2604 4272 2638
rect 4306 2604 4362 2638
rect 4396 2604 4452 2638
rect 4486 2604 4542 2638
rect 4576 2604 4632 2638
rect 4666 2604 4722 2638
rect 4756 2604 4812 2638
rect 4846 2604 4902 2638
rect 4936 2604 4992 2638
rect 5026 2604 5082 2638
rect 5116 2604 5172 2638
rect 5206 2604 5524 2638
rect 5558 2604 5614 2638
rect 5648 2604 5704 2638
rect 5738 2604 5794 2638
rect 5828 2604 5884 2638
rect 5918 2604 5974 2638
rect 6008 2604 6064 2638
rect 6098 2604 6154 2638
rect 6188 2604 6244 2638
rect 6278 2604 6334 2638
rect 6368 2604 6424 2638
rect 6458 2604 6514 2638
rect 6548 2604 6866 2638
rect 6900 2604 6956 2638
rect 6990 2604 7046 2638
rect 7080 2604 7136 2638
rect 7170 2604 7226 2638
rect 7260 2604 7316 2638
rect 7350 2604 7406 2638
rect 7440 2604 7496 2638
rect 7530 2604 7586 2638
rect 7620 2604 7676 2638
rect 7710 2604 7766 2638
rect 7800 2604 7856 2638
rect 7890 2604 8208 2638
rect 8242 2604 8298 2638
rect 8332 2604 8388 2638
rect 8422 2604 8478 2638
rect 8512 2604 8568 2638
rect 8602 2604 8658 2638
rect 8692 2604 8748 2638
rect 8782 2604 8838 2638
rect 8872 2604 8928 2638
rect 8962 2604 9018 2638
rect 9052 2604 9108 2638
rect 9142 2604 9198 2638
rect 9232 2604 9366 2638
rect 26 2483 9366 2604
rect 26 2460 156 2483
rect 26 2426 60 2460
rect 94 2449 156 2460
rect 190 2449 246 2483
rect 280 2449 336 2483
rect 370 2449 426 2483
rect 460 2449 516 2483
rect 550 2449 606 2483
rect 640 2449 696 2483
rect 730 2449 786 2483
rect 820 2449 876 2483
rect 910 2449 966 2483
rect 1000 2449 1056 2483
rect 1090 2449 1146 2483
rect 1180 2460 1498 2483
rect 1180 2449 1247 2460
rect 94 2426 1247 2449
rect 1281 2426 1402 2460
rect 1436 2449 1498 2460
rect 1532 2449 1588 2483
rect 1622 2449 1678 2483
rect 1712 2449 1768 2483
rect 1802 2449 1858 2483
rect 1892 2449 1948 2483
rect 1982 2449 2038 2483
rect 2072 2449 2128 2483
rect 2162 2449 2218 2483
rect 2252 2449 2308 2483
rect 2342 2449 2398 2483
rect 2432 2449 2488 2483
rect 2522 2460 2840 2483
rect 2522 2449 2589 2460
rect 1436 2426 2589 2449
rect 2623 2426 2744 2460
rect 2778 2449 2840 2460
rect 2874 2449 2930 2483
rect 2964 2449 3020 2483
rect 3054 2449 3110 2483
rect 3144 2449 3200 2483
rect 3234 2449 3290 2483
rect 3324 2449 3380 2483
rect 3414 2449 3470 2483
rect 3504 2449 3560 2483
rect 3594 2449 3650 2483
rect 3684 2449 3740 2483
rect 3774 2449 3830 2483
rect 3864 2460 4182 2483
rect 3864 2449 3931 2460
rect 2778 2426 3931 2449
rect 3965 2426 4086 2460
rect 4120 2449 4182 2460
rect 4216 2449 4272 2483
rect 4306 2449 4362 2483
rect 4396 2449 4452 2483
rect 4486 2449 4542 2483
rect 4576 2449 4632 2483
rect 4666 2449 4722 2483
rect 4756 2449 4812 2483
rect 4846 2449 4902 2483
rect 4936 2449 4992 2483
rect 5026 2449 5082 2483
rect 5116 2449 5172 2483
rect 5206 2460 5524 2483
rect 5206 2449 5273 2460
rect 4120 2426 5273 2449
rect 5307 2426 5428 2460
rect 5462 2449 5524 2460
rect 5558 2449 5614 2483
rect 5648 2449 5704 2483
rect 5738 2449 5794 2483
rect 5828 2449 5884 2483
rect 5918 2449 5974 2483
rect 6008 2449 6064 2483
rect 6098 2449 6154 2483
rect 6188 2449 6244 2483
rect 6278 2449 6334 2483
rect 6368 2449 6424 2483
rect 6458 2449 6514 2483
rect 6548 2460 6866 2483
rect 6548 2449 6615 2460
rect 5462 2426 6615 2449
rect 6649 2426 6770 2460
rect 6804 2449 6866 2460
rect 6900 2449 6956 2483
rect 6990 2449 7046 2483
rect 7080 2449 7136 2483
rect 7170 2449 7226 2483
rect 7260 2449 7316 2483
rect 7350 2449 7406 2483
rect 7440 2449 7496 2483
rect 7530 2449 7586 2483
rect 7620 2449 7676 2483
rect 7710 2449 7766 2483
rect 7800 2449 7856 2483
rect 7890 2460 8208 2483
rect 7890 2449 7957 2460
rect 6804 2426 7957 2449
rect 7991 2426 8112 2460
rect 8146 2449 8208 2460
rect 8242 2449 8298 2483
rect 8332 2449 8388 2483
rect 8422 2449 8478 2483
rect 8512 2449 8568 2483
rect 8602 2449 8658 2483
rect 8692 2449 8748 2483
rect 8782 2449 8838 2483
rect 8872 2449 8928 2483
rect 8962 2449 9018 2483
rect 9052 2449 9108 2483
rect 9142 2449 9198 2483
rect 9232 2460 9366 2483
rect 9232 2449 9299 2460
rect 8146 2426 9299 2449
rect 9333 2426 9366 2460
rect 26 2370 9366 2426
rect 26 2336 60 2370
rect 94 2336 1247 2370
rect 1281 2336 1402 2370
rect 1436 2336 2589 2370
rect 2623 2336 2744 2370
rect 2778 2336 3931 2370
rect 3965 2336 4086 2370
rect 4120 2336 5273 2370
rect 5307 2336 5428 2370
rect 5462 2336 6615 2370
rect 6649 2336 6770 2370
rect 6804 2336 7957 2370
rect 7991 2336 8112 2370
rect 8146 2336 9299 2370
rect 9333 2336 9366 2370
rect 26 2302 320 2336
rect 354 2302 410 2336
rect 444 2302 500 2336
rect 534 2302 590 2336
rect 624 2302 680 2336
rect 714 2302 770 2336
rect 804 2302 860 2336
rect 894 2302 950 2336
rect 984 2302 1040 2336
rect 1074 2302 1662 2336
rect 1696 2302 1752 2336
rect 1786 2302 1842 2336
rect 1876 2302 1932 2336
rect 1966 2302 2022 2336
rect 2056 2302 2112 2336
rect 2146 2302 2202 2336
rect 2236 2302 2292 2336
rect 2326 2302 2382 2336
rect 2416 2302 3004 2336
rect 3038 2302 3094 2336
rect 3128 2302 3184 2336
rect 3218 2302 3274 2336
rect 3308 2302 3364 2336
rect 3398 2302 3454 2336
rect 3488 2302 3544 2336
rect 3578 2302 3634 2336
rect 3668 2302 3724 2336
rect 3758 2302 4346 2336
rect 4380 2302 4436 2336
rect 4470 2302 4526 2336
rect 4560 2302 4616 2336
rect 4650 2302 4706 2336
rect 4740 2302 4796 2336
rect 4830 2302 4886 2336
rect 4920 2302 4976 2336
rect 5010 2302 5066 2336
rect 5100 2302 5688 2336
rect 5722 2302 5778 2336
rect 5812 2302 5868 2336
rect 5902 2302 5958 2336
rect 5992 2302 6048 2336
rect 6082 2302 6138 2336
rect 6172 2302 6228 2336
rect 6262 2302 6318 2336
rect 6352 2302 6408 2336
rect 6442 2302 7030 2336
rect 7064 2302 7120 2336
rect 7154 2302 7210 2336
rect 7244 2302 7300 2336
rect 7334 2302 7390 2336
rect 7424 2302 7480 2336
rect 7514 2302 7570 2336
rect 7604 2302 7660 2336
rect 7694 2302 7750 2336
rect 7784 2302 8372 2336
rect 8406 2302 8462 2336
rect 8496 2302 8552 2336
rect 8586 2302 8642 2336
rect 8676 2302 8732 2336
rect 8766 2302 8822 2336
rect 8856 2302 8912 2336
rect 8946 2302 9002 2336
rect 9036 2302 9092 2336
rect 9126 2302 9366 2336
rect 26 2283 9366 2302
rect 26 2280 261 2283
rect 26 2246 60 2280
rect 94 2279 261 2280
rect 94 2246 208 2279
rect 26 2245 208 2246
rect 242 2245 261 2279
rect 26 2190 261 2245
rect 1079 2280 1603 2283
rect 1079 2260 1247 2280
rect 1079 2226 1098 2260
rect 1132 2246 1247 2260
rect 1281 2246 1402 2280
rect 1436 2279 1603 2280
rect 1436 2246 1550 2279
rect 1132 2245 1550 2246
rect 1584 2245 1603 2279
rect 1132 2226 1603 2245
rect 26 2156 60 2190
rect 94 2189 261 2190
rect 94 2156 208 2189
rect 26 2155 208 2156
rect 242 2155 261 2189
rect 26 2100 261 2155
rect 26 2066 60 2100
rect 94 2099 261 2100
rect 94 2066 208 2099
rect 26 2065 208 2066
rect 242 2065 261 2099
rect 26 2010 261 2065
rect 26 1976 60 2010
rect 94 2009 261 2010
rect 94 1976 208 2009
rect 26 1975 208 1976
rect 242 1975 261 2009
rect 26 1920 261 1975
rect 26 1886 60 1920
rect 94 1919 261 1920
rect 94 1886 208 1919
rect 26 1885 208 1886
rect 242 1885 261 1919
rect 26 1830 261 1885
rect 26 1796 60 1830
rect 94 1829 261 1830
rect 94 1796 208 1829
rect 26 1795 208 1796
rect 242 1795 261 1829
rect 26 1740 261 1795
rect 26 1706 60 1740
rect 94 1739 261 1740
rect 94 1706 208 1739
rect 26 1705 208 1706
rect 242 1705 261 1739
rect 26 1650 261 1705
rect 26 1616 60 1650
rect 94 1649 261 1650
rect 94 1616 208 1649
rect 26 1615 208 1616
rect 242 1615 261 1649
rect 26 1560 261 1615
rect 26 1526 60 1560
rect 94 1559 261 1560
rect 94 1526 208 1559
rect 26 1525 208 1526
rect 242 1525 261 1559
rect 323 2162 1017 2221
rect 323 2128 384 2162
rect 418 2128 474 2162
rect 508 2128 564 2162
rect 598 2128 654 2162
rect 688 2128 744 2162
rect 778 2128 834 2162
rect 868 2128 924 2162
rect 958 2128 1017 2162
rect 323 2072 1017 2128
rect 323 2038 384 2072
rect 418 2038 474 2072
rect 508 2038 564 2072
rect 598 2038 654 2072
rect 688 2038 744 2072
rect 778 2038 834 2072
rect 868 2038 924 2072
rect 958 2038 1017 2072
rect 323 1982 1017 2038
rect 323 1948 384 1982
rect 418 1948 474 1982
rect 508 1948 564 1982
rect 598 1948 654 1982
rect 688 1948 744 1982
rect 778 1948 834 1982
rect 868 1948 924 1982
rect 958 1948 1017 1982
rect 323 1892 1017 1948
rect 323 1858 384 1892
rect 418 1858 474 1892
rect 508 1858 564 1892
rect 598 1858 654 1892
rect 688 1858 744 1892
rect 778 1858 834 1892
rect 868 1858 924 1892
rect 958 1858 1017 1892
rect 323 1802 1017 1858
rect 323 1768 384 1802
rect 418 1768 474 1802
rect 508 1768 564 1802
rect 598 1768 654 1802
rect 688 1768 744 1802
rect 778 1768 834 1802
rect 868 1768 924 1802
rect 958 1768 1017 1802
rect 323 1712 1017 1768
rect 323 1678 384 1712
rect 418 1678 474 1712
rect 508 1678 564 1712
rect 598 1678 654 1712
rect 688 1678 744 1712
rect 778 1678 834 1712
rect 868 1678 924 1712
rect 958 1678 1017 1712
rect 323 1622 1017 1678
rect 323 1588 384 1622
rect 418 1588 474 1622
rect 508 1588 564 1622
rect 598 1588 654 1622
rect 688 1588 744 1622
rect 778 1588 834 1622
rect 868 1588 924 1622
rect 958 1588 1017 1622
rect 323 1527 1017 1588
rect 1079 2190 1603 2226
rect 2421 2280 2945 2283
rect 2421 2260 2589 2280
rect 2421 2226 2440 2260
rect 2474 2246 2589 2260
rect 2623 2246 2744 2280
rect 2778 2279 2945 2280
rect 2778 2246 2892 2279
rect 2474 2245 2892 2246
rect 2926 2245 2945 2279
rect 2474 2226 2945 2245
rect 1079 2170 1247 2190
rect 1079 2136 1098 2170
rect 1132 2156 1247 2170
rect 1281 2156 1402 2190
rect 1436 2189 1603 2190
rect 1436 2156 1550 2189
rect 1132 2155 1550 2156
rect 1584 2155 1603 2189
rect 1132 2136 1603 2155
rect 1079 2100 1603 2136
rect 1079 2080 1247 2100
rect 1079 2046 1098 2080
rect 1132 2066 1247 2080
rect 1281 2066 1402 2100
rect 1436 2099 1603 2100
rect 1436 2066 1550 2099
rect 1132 2065 1550 2066
rect 1584 2065 1603 2099
rect 1132 2046 1603 2065
rect 1079 2010 1603 2046
rect 1079 1990 1247 2010
rect 1079 1956 1098 1990
rect 1132 1976 1247 1990
rect 1281 1976 1402 2010
rect 1436 2009 1603 2010
rect 1436 1976 1550 2009
rect 1132 1975 1550 1976
rect 1584 1975 1603 2009
rect 1132 1956 1603 1975
rect 1079 1920 1603 1956
rect 1079 1900 1247 1920
rect 1079 1866 1098 1900
rect 1132 1886 1247 1900
rect 1281 1886 1402 1920
rect 1436 1919 1603 1920
rect 1436 1886 1550 1919
rect 1132 1885 1550 1886
rect 1584 1885 1603 1919
rect 1132 1866 1603 1885
rect 1079 1830 1603 1866
rect 1079 1810 1247 1830
rect 1079 1776 1098 1810
rect 1132 1796 1247 1810
rect 1281 1796 1402 1830
rect 1436 1829 1603 1830
rect 1436 1796 1550 1829
rect 1132 1795 1550 1796
rect 1584 1795 1603 1829
rect 1132 1776 1603 1795
rect 1079 1740 1603 1776
rect 1079 1720 1247 1740
rect 1079 1686 1098 1720
rect 1132 1706 1247 1720
rect 1281 1706 1402 1740
rect 1436 1739 1603 1740
rect 1436 1706 1550 1739
rect 1132 1705 1550 1706
rect 1584 1705 1603 1739
rect 1132 1686 1603 1705
rect 1079 1650 1603 1686
rect 1079 1630 1247 1650
rect 1079 1596 1098 1630
rect 1132 1616 1247 1630
rect 1281 1616 1402 1650
rect 1436 1649 1603 1650
rect 1436 1616 1550 1649
rect 1132 1615 1550 1616
rect 1584 1615 1603 1649
rect 1132 1596 1603 1615
rect 1079 1560 1603 1596
rect 1079 1540 1247 1560
rect 26 1470 261 1525
rect 26 1436 60 1470
rect 94 1465 261 1470
rect 1079 1506 1098 1540
rect 1132 1526 1247 1540
rect 1281 1526 1402 1560
rect 1436 1559 1603 1560
rect 1436 1526 1550 1559
rect 1132 1525 1550 1526
rect 1584 1525 1603 1559
rect 1665 2162 2359 2221
rect 1665 2128 1726 2162
rect 1760 2128 1816 2162
rect 1850 2128 1906 2162
rect 1940 2128 1996 2162
rect 2030 2128 2086 2162
rect 2120 2128 2176 2162
rect 2210 2128 2266 2162
rect 2300 2128 2359 2162
rect 1665 2072 2359 2128
rect 1665 2038 1726 2072
rect 1760 2038 1816 2072
rect 1850 2038 1906 2072
rect 1940 2038 1996 2072
rect 2030 2038 2086 2072
rect 2120 2038 2176 2072
rect 2210 2038 2266 2072
rect 2300 2038 2359 2072
rect 1665 1982 2359 2038
rect 1665 1948 1726 1982
rect 1760 1948 1816 1982
rect 1850 1948 1906 1982
rect 1940 1948 1996 1982
rect 2030 1948 2086 1982
rect 2120 1948 2176 1982
rect 2210 1948 2266 1982
rect 2300 1948 2359 1982
rect 1665 1892 2359 1948
rect 1665 1858 1726 1892
rect 1760 1858 1816 1892
rect 1850 1858 1906 1892
rect 1940 1858 1996 1892
rect 2030 1858 2086 1892
rect 2120 1858 2176 1892
rect 2210 1858 2266 1892
rect 2300 1858 2359 1892
rect 1665 1802 2359 1858
rect 1665 1768 1726 1802
rect 1760 1768 1816 1802
rect 1850 1768 1906 1802
rect 1940 1768 1996 1802
rect 2030 1768 2086 1802
rect 2120 1768 2176 1802
rect 2210 1768 2266 1802
rect 2300 1768 2359 1802
rect 1665 1712 2359 1768
rect 1665 1678 1726 1712
rect 1760 1678 1816 1712
rect 1850 1678 1906 1712
rect 1940 1678 1996 1712
rect 2030 1678 2086 1712
rect 2120 1678 2176 1712
rect 2210 1678 2266 1712
rect 2300 1678 2359 1712
rect 1665 1622 2359 1678
rect 1665 1588 1726 1622
rect 1760 1588 1816 1622
rect 1850 1588 1906 1622
rect 1940 1588 1996 1622
rect 2030 1588 2086 1622
rect 2120 1588 2176 1622
rect 2210 1588 2266 1622
rect 2300 1588 2359 1622
rect 1665 1527 2359 1588
rect 2421 2190 2945 2226
rect 3763 2280 4287 2283
rect 3763 2260 3931 2280
rect 3763 2226 3782 2260
rect 3816 2246 3931 2260
rect 3965 2246 4086 2280
rect 4120 2279 4287 2280
rect 4120 2246 4234 2279
rect 3816 2245 4234 2246
rect 4268 2245 4287 2279
rect 3816 2226 4287 2245
rect 2421 2170 2589 2190
rect 2421 2136 2440 2170
rect 2474 2156 2589 2170
rect 2623 2156 2744 2190
rect 2778 2189 2945 2190
rect 2778 2156 2892 2189
rect 2474 2155 2892 2156
rect 2926 2155 2945 2189
rect 2474 2136 2945 2155
rect 2421 2100 2945 2136
rect 2421 2080 2589 2100
rect 2421 2046 2440 2080
rect 2474 2066 2589 2080
rect 2623 2066 2744 2100
rect 2778 2099 2945 2100
rect 2778 2066 2892 2099
rect 2474 2065 2892 2066
rect 2926 2065 2945 2099
rect 2474 2046 2945 2065
rect 2421 2010 2945 2046
rect 2421 1990 2589 2010
rect 2421 1956 2440 1990
rect 2474 1976 2589 1990
rect 2623 1976 2744 2010
rect 2778 2009 2945 2010
rect 2778 1976 2892 2009
rect 2474 1975 2892 1976
rect 2926 1975 2945 2009
rect 2474 1956 2945 1975
rect 2421 1920 2945 1956
rect 2421 1900 2589 1920
rect 2421 1866 2440 1900
rect 2474 1886 2589 1900
rect 2623 1886 2744 1920
rect 2778 1919 2945 1920
rect 2778 1886 2892 1919
rect 2474 1885 2892 1886
rect 2926 1885 2945 1919
rect 2474 1866 2945 1885
rect 2421 1830 2945 1866
rect 2421 1810 2589 1830
rect 2421 1776 2440 1810
rect 2474 1796 2589 1810
rect 2623 1796 2744 1830
rect 2778 1829 2945 1830
rect 2778 1796 2892 1829
rect 2474 1795 2892 1796
rect 2926 1795 2945 1829
rect 2474 1776 2945 1795
rect 2421 1740 2945 1776
rect 2421 1720 2589 1740
rect 2421 1686 2440 1720
rect 2474 1706 2589 1720
rect 2623 1706 2744 1740
rect 2778 1739 2945 1740
rect 2778 1706 2892 1739
rect 2474 1705 2892 1706
rect 2926 1705 2945 1739
rect 2474 1686 2945 1705
rect 2421 1650 2945 1686
rect 2421 1630 2589 1650
rect 2421 1596 2440 1630
rect 2474 1616 2589 1630
rect 2623 1616 2744 1650
rect 2778 1649 2945 1650
rect 2778 1616 2892 1649
rect 2474 1615 2892 1616
rect 2926 1615 2945 1649
rect 2474 1596 2945 1615
rect 2421 1560 2945 1596
rect 2421 1540 2589 1560
rect 1132 1506 1603 1525
rect 1079 1470 1603 1506
rect 1079 1465 1247 1470
rect 94 1446 1247 1465
rect 94 1436 286 1446
rect 26 1412 286 1436
rect 320 1412 376 1446
rect 410 1412 466 1446
rect 500 1412 556 1446
rect 590 1412 646 1446
rect 680 1412 736 1446
rect 770 1412 826 1446
rect 860 1412 916 1446
rect 950 1412 1006 1446
rect 1040 1436 1247 1446
rect 1281 1436 1402 1470
rect 1436 1465 1603 1470
rect 2421 1506 2440 1540
rect 2474 1526 2589 1540
rect 2623 1526 2744 1560
rect 2778 1559 2945 1560
rect 2778 1526 2892 1559
rect 2474 1525 2892 1526
rect 2926 1525 2945 1559
rect 3007 2162 3701 2221
rect 3007 2128 3068 2162
rect 3102 2128 3158 2162
rect 3192 2128 3248 2162
rect 3282 2128 3338 2162
rect 3372 2128 3428 2162
rect 3462 2128 3518 2162
rect 3552 2128 3608 2162
rect 3642 2128 3701 2162
rect 3007 2072 3701 2128
rect 3007 2038 3068 2072
rect 3102 2038 3158 2072
rect 3192 2038 3248 2072
rect 3282 2038 3338 2072
rect 3372 2038 3428 2072
rect 3462 2038 3518 2072
rect 3552 2038 3608 2072
rect 3642 2038 3701 2072
rect 3007 1982 3701 2038
rect 3007 1948 3068 1982
rect 3102 1948 3158 1982
rect 3192 1948 3248 1982
rect 3282 1948 3338 1982
rect 3372 1948 3428 1982
rect 3462 1948 3518 1982
rect 3552 1948 3608 1982
rect 3642 1948 3701 1982
rect 3007 1892 3701 1948
rect 3007 1858 3068 1892
rect 3102 1858 3158 1892
rect 3192 1858 3248 1892
rect 3282 1858 3338 1892
rect 3372 1858 3428 1892
rect 3462 1858 3518 1892
rect 3552 1858 3608 1892
rect 3642 1858 3701 1892
rect 3007 1802 3701 1858
rect 3007 1768 3068 1802
rect 3102 1768 3158 1802
rect 3192 1768 3248 1802
rect 3282 1768 3338 1802
rect 3372 1768 3428 1802
rect 3462 1768 3518 1802
rect 3552 1768 3608 1802
rect 3642 1768 3701 1802
rect 3007 1712 3701 1768
rect 3007 1678 3068 1712
rect 3102 1678 3158 1712
rect 3192 1678 3248 1712
rect 3282 1678 3338 1712
rect 3372 1678 3428 1712
rect 3462 1678 3518 1712
rect 3552 1678 3608 1712
rect 3642 1678 3701 1712
rect 3007 1622 3701 1678
rect 3007 1588 3068 1622
rect 3102 1588 3158 1622
rect 3192 1588 3248 1622
rect 3282 1588 3338 1622
rect 3372 1588 3428 1622
rect 3462 1588 3518 1622
rect 3552 1588 3608 1622
rect 3642 1588 3701 1622
rect 3007 1527 3701 1588
rect 3763 2190 4287 2226
rect 5105 2280 5629 2283
rect 5105 2260 5273 2280
rect 5105 2226 5124 2260
rect 5158 2246 5273 2260
rect 5307 2246 5428 2280
rect 5462 2279 5629 2280
rect 5462 2246 5576 2279
rect 5158 2245 5576 2246
rect 5610 2245 5629 2279
rect 5158 2226 5629 2245
rect 3763 2170 3931 2190
rect 3763 2136 3782 2170
rect 3816 2156 3931 2170
rect 3965 2156 4086 2190
rect 4120 2189 4287 2190
rect 4120 2156 4234 2189
rect 3816 2155 4234 2156
rect 4268 2155 4287 2189
rect 3816 2136 4287 2155
rect 3763 2100 4287 2136
rect 3763 2080 3931 2100
rect 3763 2046 3782 2080
rect 3816 2066 3931 2080
rect 3965 2066 4086 2100
rect 4120 2099 4287 2100
rect 4120 2066 4234 2099
rect 3816 2065 4234 2066
rect 4268 2065 4287 2099
rect 3816 2046 4287 2065
rect 3763 2010 4287 2046
rect 3763 1990 3931 2010
rect 3763 1956 3782 1990
rect 3816 1976 3931 1990
rect 3965 1976 4086 2010
rect 4120 2009 4287 2010
rect 4120 1976 4234 2009
rect 3816 1975 4234 1976
rect 4268 1975 4287 2009
rect 3816 1956 4287 1975
rect 3763 1920 4287 1956
rect 3763 1900 3931 1920
rect 3763 1866 3782 1900
rect 3816 1886 3931 1900
rect 3965 1886 4086 1920
rect 4120 1919 4287 1920
rect 4120 1886 4234 1919
rect 3816 1885 4234 1886
rect 4268 1885 4287 1919
rect 3816 1866 4287 1885
rect 3763 1830 4287 1866
rect 3763 1810 3931 1830
rect 3763 1776 3782 1810
rect 3816 1796 3931 1810
rect 3965 1796 4086 1830
rect 4120 1829 4287 1830
rect 4120 1796 4234 1829
rect 3816 1795 4234 1796
rect 4268 1795 4287 1829
rect 3816 1776 4287 1795
rect 3763 1740 4287 1776
rect 3763 1720 3931 1740
rect 3763 1686 3782 1720
rect 3816 1706 3931 1720
rect 3965 1706 4086 1740
rect 4120 1739 4287 1740
rect 4120 1706 4234 1739
rect 3816 1705 4234 1706
rect 4268 1705 4287 1739
rect 3816 1686 4287 1705
rect 3763 1650 4287 1686
rect 3763 1630 3931 1650
rect 3763 1596 3782 1630
rect 3816 1616 3931 1630
rect 3965 1616 4086 1650
rect 4120 1649 4287 1650
rect 4120 1616 4234 1649
rect 3816 1615 4234 1616
rect 4268 1615 4287 1649
rect 3816 1596 4287 1615
rect 3763 1560 4287 1596
rect 3763 1540 3931 1560
rect 2474 1506 2945 1525
rect 2421 1470 2945 1506
rect 2421 1465 2589 1470
rect 1436 1446 2589 1465
rect 1436 1436 1628 1446
rect 1040 1412 1628 1436
rect 1662 1412 1718 1446
rect 1752 1412 1808 1446
rect 1842 1412 1898 1446
rect 1932 1412 1988 1446
rect 2022 1412 2078 1446
rect 2112 1412 2168 1446
rect 2202 1412 2258 1446
rect 2292 1412 2348 1446
rect 2382 1436 2589 1446
rect 2623 1436 2744 1470
rect 2778 1465 2945 1470
rect 3763 1506 3782 1540
rect 3816 1526 3931 1540
rect 3965 1526 4086 1560
rect 4120 1559 4287 1560
rect 4120 1526 4234 1559
rect 3816 1525 4234 1526
rect 4268 1525 4287 1559
rect 4349 2162 5043 2221
rect 4349 2128 4410 2162
rect 4444 2128 4500 2162
rect 4534 2128 4590 2162
rect 4624 2128 4680 2162
rect 4714 2128 4770 2162
rect 4804 2128 4860 2162
rect 4894 2128 4950 2162
rect 4984 2128 5043 2162
rect 4349 2072 5043 2128
rect 4349 2038 4410 2072
rect 4444 2038 4500 2072
rect 4534 2038 4590 2072
rect 4624 2038 4680 2072
rect 4714 2038 4770 2072
rect 4804 2038 4860 2072
rect 4894 2038 4950 2072
rect 4984 2038 5043 2072
rect 4349 1982 5043 2038
rect 4349 1948 4410 1982
rect 4444 1948 4500 1982
rect 4534 1948 4590 1982
rect 4624 1948 4680 1982
rect 4714 1948 4770 1982
rect 4804 1948 4860 1982
rect 4894 1948 4950 1982
rect 4984 1948 5043 1982
rect 4349 1892 5043 1948
rect 4349 1858 4410 1892
rect 4444 1858 4500 1892
rect 4534 1858 4590 1892
rect 4624 1858 4680 1892
rect 4714 1858 4770 1892
rect 4804 1858 4860 1892
rect 4894 1858 4950 1892
rect 4984 1858 5043 1892
rect 4349 1802 5043 1858
rect 4349 1768 4410 1802
rect 4444 1768 4500 1802
rect 4534 1768 4590 1802
rect 4624 1768 4680 1802
rect 4714 1768 4770 1802
rect 4804 1768 4860 1802
rect 4894 1768 4950 1802
rect 4984 1768 5043 1802
rect 4349 1712 5043 1768
rect 4349 1678 4410 1712
rect 4444 1678 4500 1712
rect 4534 1678 4590 1712
rect 4624 1678 4680 1712
rect 4714 1678 4770 1712
rect 4804 1678 4860 1712
rect 4894 1678 4950 1712
rect 4984 1678 5043 1712
rect 4349 1622 5043 1678
rect 4349 1588 4410 1622
rect 4444 1588 4500 1622
rect 4534 1588 4590 1622
rect 4624 1588 4680 1622
rect 4714 1588 4770 1622
rect 4804 1588 4860 1622
rect 4894 1588 4950 1622
rect 4984 1588 5043 1622
rect 4349 1527 5043 1588
rect 5105 2190 5629 2226
rect 6447 2280 6971 2283
rect 6447 2260 6615 2280
rect 6447 2226 6466 2260
rect 6500 2246 6615 2260
rect 6649 2246 6770 2280
rect 6804 2279 6971 2280
rect 6804 2246 6918 2279
rect 6500 2245 6918 2246
rect 6952 2245 6971 2279
rect 6500 2226 6971 2245
rect 5105 2170 5273 2190
rect 5105 2136 5124 2170
rect 5158 2156 5273 2170
rect 5307 2156 5428 2190
rect 5462 2189 5629 2190
rect 5462 2156 5576 2189
rect 5158 2155 5576 2156
rect 5610 2155 5629 2189
rect 5158 2136 5629 2155
rect 5105 2100 5629 2136
rect 5105 2080 5273 2100
rect 5105 2046 5124 2080
rect 5158 2066 5273 2080
rect 5307 2066 5428 2100
rect 5462 2099 5629 2100
rect 5462 2066 5576 2099
rect 5158 2065 5576 2066
rect 5610 2065 5629 2099
rect 5158 2046 5629 2065
rect 5105 2010 5629 2046
rect 5105 1990 5273 2010
rect 5105 1956 5124 1990
rect 5158 1976 5273 1990
rect 5307 1976 5428 2010
rect 5462 2009 5629 2010
rect 5462 1976 5576 2009
rect 5158 1975 5576 1976
rect 5610 1975 5629 2009
rect 5158 1956 5629 1975
rect 5105 1920 5629 1956
rect 5105 1900 5273 1920
rect 5105 1866 5124 1900
rect 5158 1886 5273 1900
rect 5307 1886 5428 1920
rect 5462 1919 5629 1920
rect 5462 1886 5576 1919
rect 5158 1885 5576 1886
rect 5610 1885 5629 1919
rect 5158 1866 5629 1885
rect 5105 1830 5629 1866
rect 5105 1810 5273 1830
rect 5105 1776 5124 1810
rect 5158 1796 5273 1810
rect 5307 1796 5428 1830
rect 5462 1829 5629 1830
rect 5462 1796 5576 1829
rect 5158 1795 5576 1796
rect 5610 1795 5629 1829
rect 5158 1776 5629 1795
rect 5105 1740 5629 1776
rect 5105 1720 5273 1740
rect 5105 1686 5124 1720
rect 5158 1706 5273 1720
rect 5307 1706 5428 1740
rect 5462 1739 5629 1740
rect 5462 1706 5576 1739
rect 5158 1705 5576 1706
rect 5610 1705 5629 1739
rect 5158 1686 5629 1705
rect 5105 1650 5629 1686
rect 5105 1630 5273 1650
rect 5105 1596 5124 1630
rect 5158 1616 5273 1630
rect 5307 1616 5428 1650
rect 5462 1649 5629 1650
rect 5462 1616 5576 1649
rect 5158 1615 5576 1616
rect 5610 1615 5629 1649
rect 5158 1596 5629 1615
rect 5105 1560 5629 1596
rect 5105 1540 5273 1560
rect 3816 1506 4287 1525
rect 3763 1470 4287 1506
rect 3763 1465 3931 1470
rect 2778 1446 3931 1465
rect 2778 1436 2970 1446
rect 2382 1412 2970 1436
rect 3004 1412 3060 1446
rect 3094 1412 3150 1446
rect 3184 1412 3240 1446
rect 3274 1412 3330 1446
rect 3364 1412 3420 1446
rect 3454 1412 3510 1446
rect 3544 1412 3600 1446
rect 3634 1412 3690 1446
rect 3724 1436 3931 1446
rect 3965 1436 4086 1470
rect 4120 1465 4287 1470
rect 5105 1506 5124 1540
rect 5158 1526 5273 1540
rect 5307 1526 5428 1560
rect 5462 1559 5629 1560
rect 5462 1526 5576 1559
rect 5158 1525 5576 1526
rect 5610 1525 5629 1559
rect 5691 2162 6385 2221
rect 5691 2128 5752 2162
rect 5786 2128 5842 2162
rect 5876 2128 5932 2162
rect 5966 2128 6022 2162
rect 6056 2128 6112 2162
rect 6146 2128 6202 2162
rect 6236 2128 6292 2162
rect 6326 2128 6385 2162
rect 5691 2072 6385 2128
rect 5691 2038 5752 2072
rect 5786 2038 5842 2072
rect 5876 2038 5932 2072
rect 5966 2038 6022 2072
rect 6056 2038 6112 2072
rect 6146 2038 6202 2072
rect 6236 2038 6292 2072
rect 6326 2038 6385 2072
rect 5691 1982 6385 2038
rect 5691 1948 5752 1982
rect 5786 1948 5842 1982
rect 5876 1948 5932 1982
rect 5966 1948 6022 1982
rect 6056 1948 6112 1982
rect 6146 1948 6202 1982
rect 6236 1948 6292 1982
rect 6326 1948 6385 1982
rect 5691 1892 6385 1948
rect 5691 1858 5752 1892
rect 5786 1858 5842 1892
rect 5876 1858 5932 1892
rect 5966 1858 6022 1892
rect 6056 1858 6112 1892
rect 6146 1858 6202 1892
rect 6236 1858 6292 1892
rect 6326 1858 6385 1892
rect 5691 1802 6385 1858
rect 5691 1768 5752 1802
rect 5786 1768 5842 1802
rect 5876 1768 5932 1802
rect 5966 1768 6022 1802
rect 6056 1768 6112 1802
rect 6146 1768 6202 1802
rect 6236 1768 6292 1802
rect 6326 1768 6385 1802
rect 5691 1712 6385 1768
rect 5691 1678 5752 1712
rect 5786 1678 5842 1712
rect 5876 1678 5932 1712
rect 5966 1678 6022 1712
rect 6056 1678 6112 1712
rect 6146 1678 6202 1712
rect 6236 1678 6292 1712
rect 6326 1678 6385 1712
rect 5691 1622 6385 1678
rect 5691 1588 5752 1622
rect 5786 1588 5842 1622
rect 5876 1588 5932 1622
rect 5966 1588 6022 1622
rect 6056 1588 6112 1622
rect 6146 1588 6202 1622
rect 6236 1588 6292 1622
rect 6326 1588 6385 1622
rect 5691 1527 6385 1588
rect 6447 2190 6971 2226
rect 7789 2280 8313 2283
rect 7789 2260 7957 2280
rect 7789 2226 7808 2260
rect 7842 2246 7957 2260
rect 7991 2246 8112 2280
rect 8146 2279 8313 2280
rect 8146 2246 8260 2279
rect 7842 2245 8260 2246
rect 8294 2245 8313 2279
rect 7842 2226 8313 2245
rect 6447 2170 6615 2190
rect 6447 2136 6466 2170
rect 6500 2156 6615 2170
rect 6649 2156 6770 2190
rect 6804 2189 6971 2190
rect 6804 2156 6918 2189
rect 6500 2155 6918 2156
rect 6952 2155 6971 2189
rect 6500 2136 6971 2155
rect 6447 2100 6971 2136
rect 6447 2080 6615 2100
rect 6447 2046 6466 2080
rect 6500 2066 6615 2080
rect 6649 2066 6770 2100
rect 6804 2099 6971 2100
rect 6804 2066 6918 2099
rect 6500 2065 6918 2066
rect 6952 2065 6971 2099
rect 6500 2046 6971 2065
rect 6447 2010 6971 2046
rect 6447 1990 6615 2010
rect 6447 1956 6466 1990
rect 6500 1976 6615 1990
rect 6649 1976 6770 2010
rect 6804 2009 6971 2010
rect 6804 1976 6918 2009
rect 6500 1975 6918 1976
rect 6952 1975 6971 2009
rect 6500 1956 6971 1975
rect 6447 1920 6971 1956
rect 6447 1900 6615 1920
rect 6447 1866 6466 1900
rect 6500 1886 6615 1900
rect 6649 1886 6770 1920
rect 6804 1919 6971 1920
rect 6804 1886 6918 1919
rect 6500 1885 6918 1886
rect 6952 1885 6971 1919
rect 6500 1866 6971 1885
rect 6447 1830 6971 1866
rect 6447 1810 6615 1830
rect 6447 1776 6466 1810
rect 6500 1796 6615 1810
rect 6649 1796 6770 1830
rect 6804 1829 6971 1830
rect 6804 1796 6918 1829
rect 6500 1795 6918 1796
rect 6952 1795 6971 1829
rect 6500 1776 6971 1795
rect 6447 1740 6971 1776
rect 6447 1720 6615 1740
rect 6447 1686 6466 1720
rect 6500 1706 6615 1720
rect 6649 1706 6770 1740
rect 6804 1739 6971 1740
rect 6804 1706 6918 1739
rect 6500 1705 6918 1706
rect 6952 1705 6971 1739
rect 6500 1686 6971 1705
rect 6447 1650 6971 1686
rect 6447 1630 6615 1650
rect 6447 1596 6466 1630
rect 6500 1616 6615 1630
rect 6649 1616 6770 1650
rect 6804 1649 6971 1650
rect 6804 1616 6918 1649
rect 6500 1615 6918 1616
rect 6952 1615 6971 1649
rect 6500 1596 6971 1615
rect 6447 1560 6971 1596
rect 6447 1540 6615 1560
rect 5158 1506 5629 1525
rect 5105 1470 5629 1506
rect 5105 1465 5273 1470
rect 4120 1446 5273 1465
rect 4120 1436 4312 1446
rect 3724 1412 4312 1436
rect 4346 1412 4402 1446
rect 4436 1412 4492 1446
rect 4526 1412 4582 1446
rect 4616 1412 4672 1446
rect 4706 1412 4762 1446
rect 4796 1412 4852 1446
rect 4886 1412 4942 1446
rect 4976 1412 5032 1446
rect 5066 1436 5273 1446
rect 5307 1436 5428 1470
rect 5462 1465 5629 1470
rect 6447 1506 6466 1540
rect 6500 1526 6615 1540
rect 6649 1526 6770 1560
rect 6804 1559 6971 1560
rect 6804 1526 6918 1559
rect 6500 1525 6918 1526
rect 6952 1525 6971 1559
rect 7033 2162 7727 2221
rect 7033 2128 7094 2162
rect 7128 2128 7184 2162
rect 7218 2128 7274 2162
rect 7308 2128 7364 2162
rect 7398 2128 7454 2162
rect 7488 2128 7544 2162
rect 7578 2128 7634 2162
rect 7668 2128 7727 2162
rect 7033 2072 7727 2128
rect 7033 2038 7094 2072
rect 7128 2038 7184 2072
rect 7218 2038 7274 2072
rect 7308 2038 7364 2072
rect 7398 2038 7454 2072
rect 7488 2038 7544 2072
rect 7578 2038 7634 2072
rect 7668 2038 7727 2072
rect 7033 1982 7727 2038
rect 7033 1948 7094 1982
rect 7128 1948 7184 1982
rect 7218 1948 7274 1982
rect 7308 1948 7364 1982
rect 7398 1948 7454 1982
rect 7488 1948 7544 1982
rect 7578 1948 7634 1982
rect 7668 1948 7727 1982
rect 7033 1892 7727 1948
rect 7033 1858 7094 1892
rect 7128 1858 7184 1892
rect 7218 1858 7274 1892
rect 7308 1858 7364 1892
rect 7398 1858 7454 1892
rect 7488 1858 7544 1892
rect 7578 1858 7634 1892
rect 7668 1858 7727 1892
rect 7033 1802 7727 1858
rect 7033 1768 7094 1802
rect 7128 1768 7184 1802
rect 7218 1768 7274 1802
rect 7308 1768 7364 1802
rect 7398 1768 7454 1802
rect 7488 1768 7544 1802
rect 7578 1768 7634 1802
rect 7668 1768 7727 1802
rect 7033 1712 7727 1768
rect 7033 1678 7094 1712
rect 7128 1678 7184 1712
rect 7218 1678 7274 1712
rect 7308 1678 7364 1712
rect 7398 1678 7454 1712
rect 7488 1678 7544 1712
rect 7578 1678 7634 1712
rect 7668 1678 7727 1712
rect 7033 1622 7727 1678
rect 7033 1588 7094 1622
rect 7128 1588 7184 1622
rect 7218 1588 7274 1622
rect 7308 1588 7364 1622
rect 7398 1588 7454 1622
rect 7488 1588 7544 1622
rect 7578 1588 7634 1622
rect 7668 1588 7727 1622
rect 7033 1527 7727 1588
rect 7789 2190 8313 2226
rect 9131 2280 9366 2283
rect 9131 2260 9299 2280
rect 9131 2226 9150 2260
rect 9184 2246 9299 2260
rect 9333 2246 9366 2280
rect 9184 2226 9366 2246
rect 7789 2170 7957 2190
rect 7789 2136 7808 2170
rect 7842 2156 7957 2170
rect 7991 2156 8112 2190
rect 8146 2189 8313 2190
rect 8146 2156 8260 2189
rect 7842 2155 8260 2156
rect 8294 2155 8313 2189
rect 7842 2136 8313 2155
rect 7789 2100 8313 2136
rect 7789 2080 7957 2100
rect 7789 2046 7808 2080
rect 7842 2066 7957 2080
rect 7991 2066 8112 2100
rect 8146 2099 8313 2100
rect 8146 2066 8260 2099
rect 7842 2065 8260 2066
rect 8294 2065 8313 2099
rect 7842 2046 8313 2065
rect 7789 2010 8313 2046
rect 7789 1990 7957 2010
rect 7789 1956 7808 1990
rect 7842 1976 7957 1990
rect 7991 1976 8112 2010
rect 8146 2009 8313 2010
rect 8146 1976 8260 2009
rect 7842 1975 8260 1976
rect 8294 1975 8313 2009
rect 7842 1956 8313 1975
rect 7789 1920 8313 1956
rect 7789 1900 7957 1920
rect 7789 1866 7808 1900
rect 7842 1886 7957 1900
rect 7991 1886 8112 1920
rect 8146 1919 8313 1920
rect 8146 1886 8260 1919
rect 7842 1885 8260 1886
rect 8294 1885 8313 1919
rect 7842 1866 8313 1885
rect 7789 1830 8313 1866
rect 7789 1810 7957 1830
rect 7789 1776 7808 1810
rect 7842 1796 7957 1810
rect 7991 1796 8112 1830
rect 8146 1829 8313 1830
rect 8146 1796 8260 1829
rect 7842 1795 8260 1796
rect 8294 1795 8313 1829
rect 7842 1776 8313 1795
rect 7789 1740 8313 1776
rect 7789 1720 7957 1740
rect 7789 1686 7808 1720
rect 7842 1706 7957 1720
rect 7991 1706 8112 1740
rect 8146 1739 8313 1740
rect 8146 1706 8260 1739
rect 7842 1705 8260 1706
rect 8294 1705 8313 1739
rect 7842 1686 8313 1705
rect 7789 1650 8313 1686
rect 7789 1630 7957 1650
rect 7789 1596 7808 1630
rect 7842 1616 7957 1630
rect 7991 1616 8112 1650
rect 8146 1649 8313 1650
rect 8146 1616 8260 1649
rect 7842 1615 8260 1616
rect 8294 1615 8313 1649
rect 7842 1596 8313 1615
rect 7789 1560 8313 1596
rect 7789 1540 7957 1560
rect 6500 1506 6971 1525
rect 6447 1470 6971 1506
rect 6447 1465 6615 1470
rect 5462 1446 6615 1465
rect 5462 1436 5654 1446
rect 5066 1412 5654 1436
rect 5688 1412 5744 1446
rect 5778 1412 5834 1446
rect 5868 1412 5924 1446
rect 5958 1412 6014 1446
rect 6048 1412 6104 1446
rect 6138 1412 6194 1446
rect 6228 1412 6284 1446
rect 6318 1412 6374 1446
rect 6408 1436 6615 1446
rect 6649 1436 6770 1470
rect 6804 1465 6971 1470
rect 7789 1506 7808 1540
rect 7842 1526 7957 1540
rect 7991 1526 8112 1560
rect 8146 1559 8313 1560
rect 8146 1526 8260 1559
rect 7842 1525 8260 1526
rect 8294 1525 8313 1559
rect 8375 2162 9069 2221
rect 8375 2128 8436 2162
rect 8470 2128 8526 2162
rect 8560 2128 8616 2162
rect 8650 2128 8706 2162
rect 8740 2128 8796 2162
rect 8830 2128 8886 2162
rect 8920 2128 8976 2162
rect 9010 2128 9069 2162
rect 8375 2072 9069 2128
rect 8375 2038 8436 2072
rect 8470 2038 8526 2072
rect 8560 2038 8616 2072
rect 8650 2038 8706 2072
rect 8740 2038 8796 2072
rect 8830 2038 8886 2072
rect 8920 2038 8976 2072
rect 9010 2038 9069 2072
rect 8375 1982 9069 2038
rect 8375 1948 8436 1982
rect 8470 1948 8526 1982
rect 8560 1948 8616 1982
rect 8650 1948 8706 1982
rect 8740 1948 8796 1982
rect 8830 1948 8886 1982
rect 8920 1948 8976 1982
rect 9010 1948 9069 1982
rect 8375 1892 9069 1948
rect 8375 1858 8436 1892
rect 8470 1858 8526 1892
rect 8560 1858 8616 1892
rect 8650 1858 8706 1892
rect 8740 1858 8796 1892
rect 8830 1858 8886 1892
rect 8920 1858 8976 1892
rect 9010 1858 9069 1892
rect 8375 1802 9069 1858
rect 8375 1768 8436 1802
rect 8470 1768 8526 1802
rect 8560 1768 8616 1802
rect 8650 1768 8706 1802
rect 8740 1768 8796 1802
rect 8830 1768 8886 1802
rect 8920 1768 8976 1802
rect 9010 1768 9069 1802
rect 8375 1712 9069 1768
rect 8375 1678 8436 1712
rect 8470 1678 8526 1712
rect 8560 1678 8616 1712
rect 8650 1678 8706 1712
rect 8740 1678 8796 1712
rect 8830 1678 8886 1712
rect 8920 1678 8976 1712
rect 9010 1678 9069 1712
rect 8375 1622 9069 1678
rect 8375 1588 8436 1622
rect 8470 1588 8526 1622
rect 8560 1588 8616 1622
rect 8650 1588 8706 1622
rect 8740 1588 8796 1622
rect 8830 1588 8886 1622
rect 8920 1588 8976 1622
rect 9010 1588 9069 1622
rect 8375 1527 9069 1588
rect 9131 2190 9366 2226
rect 9131 2170 9299 2190
rect 9131 2136 9150 2170
rect 9184 2156 9299 2170
rect 9333 2156 9366 2190
rect 9184 2136 9366 2156
rect 9131 2100 9366 2136
rect 9131 2080 9299 2100
rect 9131 2046 9150 2080
rect 9184 2066 9299 2080
rect 9333 2066 9366 2100
rect 9184 2046 9366 2066
rect 9131 2010 9366 2046
rect 9131 1990 9299 2010
rect 9131 1956 9150 1990
rect 9184 1976 9299 1990
rect 9333 1976 9366 2010
rect 9184 1956 9366 1976
rect 9131 1920 9366 1956
rect 9131 1900 9299 1920
rect 9131 1866 9150 1900
rect 9184 1886 9299 1900
rect 9333 1886 9366 1920
rect 9184 1866 9366 1886
rect 9131 1830 9366 1866
rect 9131 1810 9299 1830
rect 9131 1776 9150 1810
rect 9184 1796 9299 1810
rect 9333 1796 9366 1830
rect 9184 1776 9366 1796
rect 9131 1740 9366 1776
rect 9131 1720 9299 1740
rect 9131 1686 9150 1720
rect 9184 1706 9299 1720
rect 9333 1706 9366 1740
rect 9184 1686 9366 1706
rect 9131 1650 9366 1686
rect 9131 1630 9299 1650
rect 9131 1596 9150 1630
rect 9184 1616 9299 1630
rect 9333 1616 9366 1650
rect 9184 1596 9366 1616
rect 9131 1560 9366 1596
rect 9131 1540 9299 1560
rect 7842 1506 8313 1525
rect 7789 1470 8313 1506
rect 7789 1465 7957 1470
rect 6804 1446 7957 1465
rect 6804 1436 6996 1446
rect 6408 1412 6996 1436
rect 7030 1412 7086 1446
rect 7120 1412 7176 1446
rect 7210 1412 7266 1446
rect 7300 1412 7356 1446
rect 7390 1412 7446 1446
rect 7480 1412 7536 1446
rect 7570 1412 7626 1446
rect 7660 1412 7716 1446
rect 7750 1436 7957 1446
rect 7991 1436 8112 1470
rect 8146 1465 8313 1470
rect 9131 1506 9150 1540
rect 9184 1526 9299 1540
rect 9333 1526 9366 1560
rect 9184 1506 9366 1526
rect 9131 1470 9366 1506
rect 9131 1465 9299 1470
rect 8146 1446 9299 1465
rect 8146 1436 8338 1446
rect 7750 1412 8338 1436
rect 8372 1412 8428 1446
rect 8462 1412 8518 1446
rect 8552 1412 8608 1446
rect 8642 1412 8698 1446
rect 8732 1412 8788 1446
rect 8822 1412 8878 1446
rect 8912 1412 8968 1446
rect 9002 1412 9058 1446
rect 9092 1436 9299 1446
rect 9333 1436 9366 1470
rect 9092 1412 9366 1436
rect 26 1380 9366 1412
rect 26 1346 60 1380
rect 94 1346 1247 1380
rect 1281 1346 1402 1380
rect 1436 1346 2589 1380
rect 2623 1346 2744 1380
rect 2778 1346 3931 1380
rect 3965 1346 4086 1380
rect 4120 1346 5273 1380
rect 5307 1346 5428 1380
rect 5462 1346 6615 1380
rect 6649 1346 6770 1380
rect 6804 1346 7957 1380
rect 7991 1346 8112 1380
rect 8146 1346 9299 1380
rect 9333 1346 9366 1380
rect 26 1296 9366 1346
rect 26 1262 156 1296
rect 190 1262 246 1296
rect 280 1262 336 1296
rect 370 1262 426 1296
rect 460 1262 516 1296
rect 550 1262 606 1296
rect 640 1262 696 1296
rect 730 1262 786 1296
rect 820 1262 876 1296
rect 910 1262 966 1296
rect 1000 1262 1056 1296
rect 1090 1262 1146 1296
rect 1180 1262 1498 1296
rect 1532 1262 1588 1296
rect 1622 1262 1678 1296
rect 1712 1262 1768 1296
rect 1802 1262 1858 1296
rect 1892 1262 1948 1296
rect 1982 1262 2038 1296
rect 2072 1262 2128 1296
rect 2162 1262 2218 1296
rect 2252 1262 2308 1296
rect 2342 1262 2398 1296
rect 2432 1262 2488 1296
rect 2522 1262 2840 1296
rect 2874 1262 2930 1296
rect 2964 1262 3020 1296
rect 3054 1262 3110 1296
rect 3144 1262 3200 1296
rect 3234 1262 3290 1296
rect 3324 1262 3380 1296
rect 3414 1262 3470 1296
rect 3504 1262 3560 1296
rect 3594 1262 3650 1296
rect 3684 1262 3740 1296
rect 3774 1262 3830 1296
rect 3864 1262 4182 1296
rect 4216 1262 4272 1296
rect 4306 1262 4362 1296
rect 4396 1262 4452 1296
rect 4486 1262 4542 1296
rect 4576 1262 4632 1296
rect 4666 1262 4722 1296
rect 4756 1262 4812 1296
rect 4846 1262 4902 1296
rect 4936 1262 4992 1296
rect 5026 1262 5082 1296
rect 5116 1262 5172 1296
rect 5206 1262 5524 1296
rect 5558 1262 5614 1296
rect 5648 1262 5704 1296
rect 5738 1262 5794 1296
rect 5828 1262 5884 1296
rect 5918 1262 5974 1296
rect 6008 1262 6064 1296
rect 6098 1262 6154 1296
rect 6188 1262 6244 1296
rect 6278 1262 6334 1296
rect 6368 1262 6424 1296
rect 6458 1262 6514 1296
rect 6548 1262 6866 1296
rect 6900 1262 6956 1296
rect 6990 1262 7046 1296
rect 7080 1262 7136 1296
rect 7170 1262 7226 1296
rect 7260 1262 7316 1296
rect 7350 1262 7406 1296
rect 7440 1262 7496 1296
rect 7530 1262 7586 1296
rect 7620 1262 7676 1296
rect 7710 1262 7766 1296
rect 7800 1262 7856 1296
rect 7890 1262 8208 1296
rect 8242 1262 8298 1296
rect 8332 1262 8388 1296
rect 8422 1262 8478 1296
rect 8512 1262 8568 1296
rect 8602 1262 8658 1296
rect 8692 1262 8748 1296
rect 8782 1262 8838 1296
rect 8872 1262 8928 1296
rect 8962 1262 9018 1296
rect 9052 1262 9108 1296
rect 9142 1262 9198 1296
rect 9232 1262 9366 1296
rect 26 1141 9366 1262
rect 26 1118 6866 1141
rect 26 1084 6770 1118
rect 6804 1107 6866 1118
rect 6900 1107 6956 1141
rect 6990 1107 7046 1141
rect 7080 1107 7136 1141
rect 7170 1107 7226 1141
rect 7260 1107 7316 1141
rect 7350 1107 7406 1141
rect 7440 1107 7496 1141
rect 7530 1107 7586 1141
rect 7620 1107 7676 1141
rect 7710 1107 7766 1141
rect 7800 1107 7856 1141
rect 7890 1118 8208 1141
rect 7890 1107 7957 1118
rect 6804 1084 7957 1107
rect 7991 1084 8112 1118
rect 8146 1107 8208 1118
rect 8242 1107 8298 1141
rect 8332 1107 8388 1141
rect 8422 1107 8478 1141
rect 8512 1107 8568 1141
rect 8602 1107 8658 1141
rect 8692 1107 8748 1141
rect 8782 1107 8838 1141
rect 8872 1107 8928 1141
rect 8962 1107 9018 1141
rect 9052 1107 9108 1141
rect 9142 1107 9198 1141
rect 9232 1118 9366 1141
rect 9232 1107 9299 1118
rect 8146 1084 9299 1107
rect 9333 1084 9366 1118
rect 26 1028 9366 1084
rect 26 994 6770 1028
rect 6804 994 7957 1028
rect 7991 994 8112 1028
rect 8146 994 9299 1028
rect 9333 994 9366 1028
rect 26 960 7030 994
rect 7064 960 7120 994
rect 7154 960 7210 994
rect 7244 960 7300 994
rect 7334 960 7390 994
rect 7424 960 7480 994
rect 7514 960 7570 994
rect 7604 960 7660 994
rect 7694 960 7750 994
rect 7784 960 8372 994
rect 8406 960 8462 994
rect 8496 960 8552 994
rect 8586 960 8642 994
rect 8676 960 8732 994
rect 8766 960 8822 994
rect 8856 960 8912 994
rect 8946 960 9002 994
rect 9036 960 9092 994
rect 9126 960 9366 994
rect 26 941 9366 960
rect 26 123 261 941
rect 1079 123 1603 941
rect 2421 123 2945 941
rect 3763 123 4287 941
rect 5105 123 5629 941
rect 6447 938 6971 941
rect 6447 904 6770 938
rect 6804 937 6971 938
rect 6804 904 6918 937
rect 6447 903 6918 904
rect 6952 903 6971 937
rect 6447 848 6971 903
rect 7789 938 8313 941
rect 7789 918 7957 938
rect 7789 884 7808 918
rect 7842 904 7957 918
rect 7991 904 8112 938
rect 8146 937 8313 938
rect 8146 904 8260 937
rect 7842 903 8260 904
rect 8294 903 8313 937
rect 7842 884 8313 903
rect 6447 814 6770 848
rect 6804 847 6971 848
rect 6804 814 6918 847
rect 6447 813 6918 814
rect 6952 813 6971 847
rect 6447 758 6971 813
rect 6447 724 6770 758
rect 6804 757 6971 758
rect 6804 724 6918 757
rect 6447 723 6918 724
rect 6952 723 6971 757
rect 6447 668 6971 723
rect 6447 634 6770 668
rect 6804 667 6971 668
rect 6804 634 6918 667
rect 6447 633 6918 634
rect 6952 633 6971 667
rect 6447 578 6971 633
rect 6447 544 6770 578
rect 6804 577 6971 578
rect 6804 544 6918 577
rect 6447 543 6918 544
rect 6952 543 6971 577
rect 6447 488 6971 543
rect 6447 454 6770 488
rect 6804 487 6971 488
rect 6804 454 6918 487
rect 6447 453 6918 454
rect 6952 453 6971 487
rect 6447 398 6971 453
rect 6447 364 6770 398
rect 6804 397 6971 398
rect 6804 364 6918 397
rect 6447 363 6918 364
rect 6952 363 6971 397
rect 6447 308 6971 363
rect 6447 274 6770 308
rect 6804 307 6971 308
rect 6804 274 6918 307
rect 6447 273 6918 274
rect 6952 273 6971 307
rect 6447 218 6971 273
rect 6447 184 6770 218
rect 6804 217 6971 218
rect 6804 184 6918 217
rect 6447 183 6918 184
rect 6952 183 6971 217
rect 7033 820 7727 879
rect 7033 786 7094 820
rect 7128 786 7184 820
rect 7218 786 7274 820
rect 7308 786 7364 820
rect 7398 786 7454 820
rect 7488 786 7544 820
rect 7578 786 7634 820
rect 7668 786 7727 820
rect 7033 730 7727 786
rect 7033 696 7094 730
rect 7128 696 7184 730
rect 7218 696 7274 730
rect 7308 696 7364 730
rect 7398 696 7454 730
rect 7488 696 7544 730
rect 7578 696 7634 730
rect 7668 696 7727 730
rect 7033 640 7727 696
rect 7033 606 7094 640
rect 7128 606 7184 640
rect 7218 606 7274 640
rect 7308 606 7364 640
rect 7398 606 7454 640
rect 7488 606 7544 640
rect 7578 606 7634 640
rect 7668 606 7727 640
rect 7033 550 7727 606
rect 7033 516 7094 550
rect 7128 516 7184 550
rect 7218 516 7274 550
rect 7308 516 7364 550
rect 7398 516 7454 550
rect 7488 516 7544 550
rect 7578 516 7634 550
rect 7668 516 7727 550
rect 7033 460 7727 516
rect 7033 426 7094 460
rect 7128 426 7184 460
rect 7218 426 7274 460
rect 7308 426 7364 460
rect 7398 426 7454 460
rect 7488 426 7544 460
rect 7578 426 7634 460
rect 7668 426 7727 460
rect 7033 370 7727 426
rect 7033 336 7094 370
rect 7128 336 7184 370
rect 7218 336 7274 370
rect 7308 336 7364 370
rect 7398 336 7454 370
rect 7488 336 7544 370
rect 7578 336 7634 370
rect 7668 336 7727 370
rect 7033 280 7727 336
rect 7033 246 7094 280
rect 7128 246 7184 280
rect 7218 246 7274 280
rect 7308 246 7364 280
rect 7398 246 7454 280
rect 7488 246 7544 280
rect 7578 246 7634 280
rect 7668 246 7727 280
rect 7033 185 7727 246
rect 7789 848 8313 884
rect 9131 938 9366 941
rect 9131 918 9299 938
rect 9131 884 9150 918
rect 9184 904 9299 918
rect 9333 904 9366 938
rect 9184 884 9366 904
rect 7789 828 7957 848
rect 7789 794 7808 828
rect 7842 814 7957 828
rect 7991 814 8112 848
rect 8146 847 8313 848
rect 8146 814 8260 847
rect 7842 813 8260 814
rect 8294 813 8313 847
rect 7842 794 8313 813
rect 7789 758 8313 794
rect 7789 738 7957 758
rect 7789 704 7808 738
rect 7842 724 7957 738
rect 7991 724 8112 758
rect 8146 757 8313 758
rect 8146 724 8260 757
rect 7842 723 8260 724
rect 8294 723 8313 757
rect 7842 704 8313 723
rect 7789 668 8313 704
rect 7789 648 7957 668
rect 7789 614 7808 648
rect 7842 634 7957 648
rect 7991 634 8112 668
rect 8146 667 8313 668
rect 8146 634 8260 667
rect 7842 633 8260 634
rect 8294 633 8313 667
rect 7842 614 8313 633
rect 7789 578 8313 614
rect 7789 558 7957 578
rect 7789 524 7808 558
rect 7842 544 7957 558
rect 7991 544 8112 578
rect 8146 577 8313 578
rect 8146 544 8260 577
rect 7842 543 8260 544
rect 8294 543 8313 577
rect 7842 524 8313 543
rect 7789 488 8313 524
rect 7789 468 7957 488
rect 7789 434 7808 468
rect 7842 454 7957 468
rect 7991 454 8112 488
rect 8146 487 8313 488
rect 8146 454 8260 487
rect 7842 453 8260 454
rect 8294 453 8313 487
rect 7842 434 8313 453
rect 7789 398 8313 434
rect 7789 378 7957 398
rect 7789 344 7808 378
rect 7842 364 7957 378
rect 7991 364 8112 398
rect 8146 397 8313 398
rect 8146 364 8260 397
rect 7842 363 8260 364
rect 8294 363 8313 397
rect 7842 344 8313 363
rect 7789 308 8313 344
rect 7789 288 7957 308
rect 7789 254 7808 288
rect 7842 274 7957 288
rect 7991 274 8112 308
rect 8146 307 8313 308
rect 8146 274 8260 307
rect 7842 273 8260 274
rect 8294 273 8313 307
rect 7842 254 8313 273
rect 7789 218 8313 254
rect 7789 198 7957 218
rect 6447 128 6971 183
rect 6447 123 6770 128
rect 26 94 6770 123
rect 6804 123 6971 128
rect 7789 164 7808 198
rect 7842 184 7957 198
rect 7991 184 8112 218
rect 8146 217 8313 218
rect 8146 184 8260 217
rect 7842 183 8260 184
rect 8294 183 8313 217
rect 8375 820 9069 879
rect 8375 786 8436 820
rect 8470 786 8526 820
rect 8560 786 8616 820
rect 8650 786 8706 820
rect 8740 786 8796 820
rect 8830 786 8886 820
rect 8920 786 8976 820
rect 9010 786 9069 820
rect 8375 730 9069 786
rect 8375 696 8436 730
rect 8470 696 8526 730
rect 8560 696 8616 730
rect 8650 696 8706 730
rect 8740 696 8796 730
rect 8830 696 8886 730
rect 8920 696 8976 730
rect 9010 696 9069 730
rect 8375 640 9069 696
rect 8375 606 8436 640
rect 8470 606 8526 640
rect 8560 606 8616 640
rect 8650 606 8706 640
rect 8740 606 8796 640
rect 8830 606 8886 640
rect 8920 606 8976 640
rect 9010 606 9069 640
rect 8375 550 9069 606
rect 8375 516 8436 550
rect 8470 516 8526 550
rect 8560 516 8616 550
rect 8650 516 8706 550
rect 8740 516 8796 550
rect 8830 516 8886 550
rect 8920 516 8976 550
rect 9010 516 9069 550
rect 8375 460 9069 516
rect 8375 426 8436 460
rect 8470 426 8526 460
rect 8560 426 8616 460
rect 8650 426 8706 460
rect 8740 426 8796 460
rect 8830 426 8886 460
rect 8920 426 8976 460
rect 9010 426 9069 460
rect 8375 370 9069 426
rect 8375 336 8436 370
rect 8470 336 8526 370
rect 8560 336 8616 370
rect 8650 336 8706 370
rect 8740 336 8796 370
rect 8830 336 8886 370
rect 8920 336 8976 370
rect 9010 336 9069 370
rect 8375 280 9069 336
rect 8375 246 8436 280
rect 8470 246 8526 280
rect 8560 246 8616 280
rect 8650 246 8706 280
rect 8740 246 8796 280
rect 8830 246 8886 280
rect 8920 246 8976 280
rect 9010 246 9069 280
rect 8375 185 9069 246
rect 9131 848 9366 884
rect 9131 828 9299 848
rect 9131 794 9150 828
rect 9184 814 9299 828
rect 9333 814 9366 848
rect 9184 794 9366 814
rect 9131 758 9366 794
rect 9131 738 9299 758
rect 9131 704 9150 738
rect 9184 724 9299 738
rect 9333 724 9366 758
rect 9184 704 9366 724
rect 9131 668 9366 704
rect 9131 648 9299 668
rect 9131 614 9150 648
rect 9184 634 9299 648
rect 9333 634 9366 668
rect 9184 614 9366 634
rect 9131 578 9366 614
rect 9131 558 9299 578
rect 9131 524 9150 558
rect 9184 544 9299 558
rect 9333 544 9366 578
rect 9184 524 9366 544
rect 9131 488 9366 524
rect 9131 468 9299 488
rect 9131 434 9150 468
rect 9184 454 9299 468
rect 9333 454 9366 488
rect 9184 434 9366 454
rect 9131 398 9366 434
rect 9131 378 9299 398
rect 9131 344 9150 378
rect 9184 364 9299 378
rect 9333 364 9366 398
rect 9184 344 9366 364
rect 9131 308 9366 344
rect 9131 288 9299 308
rect 9131 254 9150 288
rect 9184 274 9299 288
rect 9333 274 9366 308
rect 9184 254 9366 274
rect 9131 218 9366 254
rect 9131 198 9299 218
rect 7842 164 8313 183
rect 7789 128 8313 164
rect 7789 123 7957 128
rect 6804 104 7957 123
rect 6804 94 6996 104
rect 26 70 6996 94
rect 7030 70 7086 104
rect 7120 70 7176 104
rect 7210 70 7266 104
rect 7300 70 7356 104
rect 7390 70 7446 104
rect 7480 70 7536 104
rect 7570 70 7626 104
rect 7660 70 7716 104
rect 7750 94 7957 104
rect 7991 94 8112 128
rect 8146 123 8313 128
rect 9131 164 9150 198
rect 9184 184 9299 198
rect 9333 184 9366 218
rect 9184 164 9366 184
rect 9131 128 9366 164
rect 9131 123 9299 128
rect 8146 104 9299 123
rect 8146 94 8338 104
rect 7750 70 8338 94
rect 8372 70 8428 104
rect 8462 70 8518 104
rect 8552 70 8608 104
rect 8642 70 8698 104
rect 8732 70 8788 104
rect 8822 70 8878 104
rect 8912 70 8968 104
rect 9002 70 9058 104
rect 9092 94 9299 104
rect 9333 94 9366 128
rect 9092 70 9366 94
rect 26 38 9366 70
rect 26 4 6770 38
rect 6804 4 7957 38
rect 7991 4 8112 38
rect 8146 4 9299 38
rect 9333 4 9366 38
rect 26 -46 9366 4
rect 26 -80 6866 -46
rect 6900 -80 6956 -46
rect 6990 -80 7046 -46
rect 7080 -80 7136 -46
rect 7170 -80 7226 -46
rect 7260 -80 7316 -46
rect 7350 -80 7406 -46
rect 7440 -80 7496 -46
rect 7530 -80 7586 -46
rect 7620 -80 7676 -46
rect 7710 -80 7766 -46
rect 7800 -80 7856 -46
rect 7890 -80 8208 -46
rect 8242 -80 8298 -46
rect 8332 -80 8388 -46
rect 8422 -80 8478 -46
rect 8512 -80 8568 -46
rect 8602 -80 8658 -46
rect 8692 -80 8748 -46
rect 8782 -80 8838 -46
rect 8872 -80 8928 -46
rect 8962 -80 9018 -46
rect 9052 -80 9108 -46
rect 9142 -80 9198 -46
rect 9232 -80 9366 -46
rect 26 -201 9366 -80
rect 26 -224 6866 -201
rect 26 -258 6770 -224
rect 6804 -235 6866 -224
rect 6900 -235 6956 -201
rect 6990 -235 7046 -201
rect 7080 -235 7136 -201
rect 7170 -235 7226 -201
rect 7260 -235 7316 -201
rect 7350 -235 7406 -201
rect 7440 -235 7496 -201
rect 7530 -235 7586 -201
rect 7620 -235 7676 -201
rect 7710 -235 7766 -201
rect 7800 -235 7856 -201
rect 7890 -224 8208 -201
rect 7890 -235 7957 -224
rect 6804 -258 7957 -235
rect 7991 -258 8112 -224
rect 8146 -235 8208 -224
rect 8242 -235 8298 -201
rect 8332 -235 8388 -201
rect 8422 -235 8478 -201
rect 8512 -235 8568 -201
rect 8602 -235 8658 -201
rect 8692 -235 8748 -201
rect 8782 -235 8838 -201
rect 8872 -235 8928 -201
rect 8962 -235 9018 -201
rect 9052 -235 9108 -201
rect 9142 -235 9198 -201
rect 9232 -224 9366 -201
rect 9232 -235 9299 -224
rect 8146 -258 9299 -235
rect 9333 -258 9366 -224
rect 26 -314 9366 -258
rect 26 -348 6770 -314
rect 6804 -348 7957 -314
rect 7991 -348 8112 -314
rect 8146 -348 9299 -314
rect 9333 -348 9366 -314
rect 26 -382 7030 -348
rect 7064 -382 7120 -348
rect 7154 -382 7210 -348
rect 7244 -382 7300 -348
rect 7334 -382 7390 -348
rect 7424 -382 7480 -348
rect 7514 -382 7570 -348
rect 7604 -382 7660 -348
rect 7694 -382 7750 -348
rect 7784 -382 8372 -348
rect 8406 -382 8462 -348
rect 8496 -382 8552 -348
rect 8586 -382 8642 -348
rect 8676 -382 8732 -348
rect 8766 -382 8822 -348
rect 8856 -382 8912 -348
rect 8946 -382 9002 -348
rect 9036 -382 9092 -348
rect 9126 -382 9366 -348
rect 26 -401 9366 -382
rect 26 -1219 261 -401
rect 1079 -1219 1603 -401
rect 2421 -1219 2945 -401
rect 3763 -1219 4287 -401
rect 5105 -1219 5629 -401
rect 6447 -404 6971 -401
rect 6447 -438 6770 -404
rect 6804 -405 6971 -404
rect 6804 -438 6918 -405
rect 6447 -439 6918 -438
rect 6952 -439 6971 -405
rect 6447 -494 6971 -439
rect 7789 -404 8313 -401
rect 7789 -424 7957 -404
rect 7789 -458 7808 -424
rect 7842 -438 7957 -424
rect 7991 -438 8112 -404
rect 8146 -405 8313 -404
rect 8146 -438 8260 -405
rect 7842 -439 8260 -438
rect 8294 -439 8313 -405
rect 7842 -458 8313 -439
rect 6447 -528 6770 -494
rect 6804 -495 6971 -494
rect 6804 -528 6918 -495
rect 6447 -529 6918 -528
rect 6952 -529 6971 -495
rect 6447 -584 6971 -529
rect 6447 -618 6770 -584
rect 6804 -585 6971 -584
rect 6804 -618 6918 -585
rect 6447 -619 6918 -618
rect 6952 -619 6971 -585
rect 6447 -674 6971 -619
rect 6447 -708 6770 -674
rect 6804 -675 6971 -674
rect 6804 -708 6918 -675
rect 6447 -709 6918 -708
rect 6952 -709 6971 -675
rect 6447 -764 6971 -709
rect 6447 -798 6770 -764
rect 6804 -765 6971 -764
rect 6804 -798 6918 -765
rect 6447 -799 6918 -798
rect 6952 -799 6971 -765
rect 6447 -854 6971 -799
rect 6447 -888 6770 -854
rect 6804 -855 6971 -854
rect 6804 -888 6918 -855
rect 6447 -889 6918 -888
rect 6952 -889 6971 -855
rect 6447 -944 6971 -889
rect 6447 -978 6770 -944
rect 6804 -945 6971 -944
rect 6804 -978 6918 -945
rect 6447 -979 6918 -978
rect 6952 -979 6971 -945
rect 6447 -1034 6971 -979
rect 6447 -1068 6770 -1034
rect 6804 -1035 6971 -1034
rect 6804 -1068 6918 -1035
rect 6447 -1069 6918 -1068
rect 6952 -1069 6971 -1035
rect 6447 -1124 6971 -1069
rect 6447 -1158 6770 -1124
rect 6804 -1125 6971 -1124
rect 6804 -1158 6918 -1125
rect 6447 -1159 6918 -1158
rect 6952 -1159 6971 -1125
rect 7033 -522 7727 -463
rect 7033 -556 7094 -522
rect 7128 -556 7184 -522
rect 7218 -556 7274 -522
rect 7308 -556 7364 -522
rect 7398 -556 7454 -522
rect 7488 -556 7544 -522
rect 7578 -556 7634 -522
rect 7668 -556 7727 -522
rect 7033 -612 7727 -556
rect 7033 -646 7094 -612
rect 7128 -646 7184 -612
rect 7218 -646 7274 -612
rect 7308 -646 7364 -612
rect 7398 -646 7454 -612
rect 7488 -646 7544 -612
rect 7578 -646 7634 -612
rect 7668 -646 7727 -612
rect 7033 -702 7727 -646
rect 7033 -736 7094 -702
rect 7128 -736 7184 -702
rect 7218 -736 7274 -702
rect 7308 -736 7364 -702
rect 7398 -736 7454 -702
rect 7488 -736 7544 -702
rect 7578 -736 7634 -702
rect 7668 -736 7727 -702
rect 7033 -792 7727 -736
rect 7033 -826 7094 -792
rect 7128 -826 7184 -792
rect 7218 -826 7274 -792
rect 7308 -826 7364 -792
rect 7398 -826 7454 -792
rect 7488 -826 7544 -792
rect 7578 -826 7634 -792
rect 7668 -826 7727 -792
rect 7033 -882 7727 -826
rect 7033 -916 7094 -882
rect 7128 -916 7184 -882
rect 7218 -916 7274 -882
rect 7308 -916 7364 -882
rect 7398 -916 7454 -882
rect 7488 -916 7544 -882
rect 7578 -916 7634 -882
rect 7668 -916 7727 -882
rect 7033 -972 7727 -916
rect 7033 -1006 7094 -972
rect 7128 -1006 7184 -972
rect 7218 -1006 7274 -972
rect 7308 -1006 7364 -972
rect 7398 -1006 7454 -972
rect 7488 -1006 7544 -972
rect 7578 -1006 7634 -972
rect 7668 -1006 7727 -972
rect 7033 -1062 7727 -1006
rect 7033 -1096 7094 -1062
rect 7128 -1096 7184 -1062
rect 7218 -1096 7274 -1062
rect 7308 -1096 7364 -1062
rect 7398 -1096 7454 -1062
rect 7488 -1096 7544 -1062
rect 7578 -1096 7634 -1062
rect 7668 -1096 7727 -1062
rect 7033 -1157 7727 -1096
rect 7789 -494 8313 -458
rect 9131 -404 9366 -401
rect 9131 -424 9299 -404
rect 9131 -458 9150 -424
rect 9184 -438 9299 -424
rect 9333 -438 9366 -404
rect 9184 -458 9366 -438
rect 7789 -514 7957 -494
rect 7789 -548 7808 -514
rect 7842 -528 7957 -514
rect 7991 -528 8112 -494
rect 8146 -495 8313 -494
rect 8146 -528 8260 -495
rect 7842 -529 8260 -528
rect 8294 -529 8313 -495
rect 7842 -548 8313 -529
rect 7789 -584 8313 -548
rect 7789 -604 7957 -584
rect 7789 -638 7808 -604
rect 7842 -618 7957 -604
rect 7991 -618 8112 -584
rect 8146 -585 8313 -584
rect 8146 -618 8260 -585
rect 7842 -619 8260 -618
rect 8294 -619 8313 -585
rect 7842 -638 8313 -619
rect 7789 -674 8313 -638
rect 7789 -694 7957 -674
rect 7789 -728 7808 -694
rect 7842 -708 7957 -694
rect 7991 -708 8112 -674
rect 8146 -675 8313 -674
rect 8146 -708 8260 -675
rect 7842 -709 8260 -708
rect 8294 -709 8313 -675
rect 7842 -728 8313 -709
rect 7789 -764 8313 -728
rect 7789 -784 7957 -764
rect 7789 -818 7808 -784
rect 7842 -798 7957 -784
rect 7991 -798 8112 -764
rect 8146 -765 8313 -764
rect 8146 -798 8260 -765
rect 7842 -799 8260 -798
rect 8294 -799 8313 -765
rect 7842 -818 8313 -799
rect 7789 -854 8313 -818
rect 7789 -874 7957 -854
rect 7789 -908 7808 -874
rect 7842 -888 7957 -874
rect 7991 -888 8112 -854
rect 8146 -855 8313 -854
rect 8146 -888 8260 -855
rect 7842 -889 8260 -888
rect 8294 -889 8313 -855
rect 7842 -908 8313 -889
rect 7789 -944 8313 -908
rect 7789 -964 7957 -944
rect 7789 -998 7808 -964
rect 7842 -978 7957 -964
rect 7991 -978 8112 -944
rect 8146 -945 8313 -944
rect 8146 -978 8260 -945
rect 7842 -979 8260 -978
rect 8294 -979 8313 -945
rect 7842 -998 8313 -979
rect 7789 -1034 8313 -998
rect 7789 -1054 7957 -1034
rect 7789 -1088 7808 -1054
rect 7842 -1068 7957 -1054
rect 7991 -1068 8112 -1034
rect 8146 -1035 8313 -1034
rect 8146 -1068 8260 -1035
rect 7842 -1069 8260 -1068
rect 8294 -1069 8313 -1035
rect 7842 -1088 8313 -1069
rect 7789 -1124 8313 -1088
rect 7789 -1144 7957 -1124
rect 6447 -1214 6971 -1159
rect 6447 -1219 6770 -1214
rect 26 -1248 6770 -1219
rect 6804 -1219 6971 -1214
rect 7789 -1178 7808 -1144
rect 7842 -1158 7957 -1144
rect 7991 -1158 8112 -1124
rect 8146 -1125 8313 -1124
rect 8146 -1158 8260 -1125
rect 7842 -1159 8260 -1158
rect 8294 -1159 8313 -1125
rect 8375 -522 9069 -463
rect 8375 -556 8436 -522
rect 8470 -556 8526 -522
rect 8560 -556 8616 -522
rect 8650 -556 8706 -522
rect 8740 -556 8796 -522
rect 8830 -556 8886 -522
rect 8920 -556 8976 -522
rect 9010 -556 9069 -522
rect 8375 -612 9069 -556
rect 8375 -646 8436 -612
rect 8470 -646 8526 -612
rect 8560 -646 8616 -612
rect 8650 -646 8706 -612
rect 8740 -646 8796 -612
rect 8830 -646 8886 -612
rect 8920 -646 8976 -612
rect 9010 -646 9069 -612
rect 8375 -702 9069 -646
rect 8375 -736 8436 -702
rect 8470 -736 8526 -702
rect 8560 -736 8616 -702
rect 8650 -736 8706 -702
rect 8740 -736 8796 -702
rect 8830 -736 8886 -702
rect 8920 -736 8976 -702
rect 9010 -736 9069 -702
rect 8375 -792 9069 -736
rect 8375 -826 8436 -792
rect 8470 -826 8526 -792
rect 8560 -826 8616 -792
rect 8650 -826 8706 -792
rect 8740 -826 8796 -792
rect 8830 -826 8886 -792
rect 8920 -826 8976 -792
rect 9010 -826 9069 -792
rect 8375 -882 9069 -826
rect 8375 -916 8436 -882
rect 8470 -916 8526 -882
rect 8560 -916 8616 -882
rect 8650 -916 8706 -882
rect 8740 -916 8796 -882
rect 8830 -916 8886 -882
rect 8920 -916 8976 -882
rect 9010 -916 9069 -882
rect 8375 -972 9069 -916
rect 8375 -1006 8436 -972
rect 8470 -1006 8526 -972
rect 8560 -1006 8616 -972
rect 8650 -1006 8706 -972
rect 8740 -1006 8796 -972
rect 8830 -1006 8886 -972
rect 8920 -1006 8976 -972
rect 9010 -1006 9069 -972
rect 8375 -1062 9069 -1006
rect 8375 -1096 8436 -1062
rect 8470 -1096 8526 -1062
rect 8560 -1096 8616 -1062
rect 8650 -1096 8706 -1062
rect 8740 -1096 8796 -1062
rect 8830 -1096 8886 -1062
rect 8920 -1096 8976 -1062
rect 9010 -1096 9069 -1062
rect 8375 -1157 9069 -1096
rect 9131 -494 9366 -458
rect 9131 -514 9299 -494
rect 9131 -548 9150 -514
rect 9184 -528 9299 -514
rect 9333 -528 9366 -494
rect 9184 -548 9366 -528
rect 9131 -584 9366 -548
rect 9131 -604 9299 -584
rect 9131 -638 9150 -604
rect 9184 -618 9299 -604
rect 9333 -618 9366 -584
rect 9184 -638 9366 -618
rect 9131 -674 9366 -638
rect 9131 -694 9299 -674
rect 9131 -728 9150 -694
rect 9184 -708 9299 -694
rect 9333 -708 9366 -674
rect 9184 -728 9366 -708
rect 9131 -764 9366 -728
rect 9131 -784 9299 -764
rect 9131 -818 9150 -784
rect 9184 -798 9299 -784
rect 9333 -798 9366 -764
rect 9184 -818 9366 -798
rect 9131 -854 9366 -818
rect 9131 -874 9299 -854
rect 9131 -908 9150 -874
rect 9184 -888 9299 -874
rect 9333 -888 9366 -854
rect 9184 -908 9366 -888
rect 9131 -944 9366 -908
rect 9131 -964 9299 -944
rect 9131 -998 9150 -964
rect 9184 -978 9299 -964
rect 9333 -978 9366 -944
rect 9184 -998 9366 -978
rect 9131 -1034 9366 -998
rect 9131 -1054 9299 -1034
rect 9131 -1088 9150 -1054
rect 9184 -1068 9299 -1054
rect 9333 -1068 9366 -1034
rect 9184 -1088 9366 -1068
rect 9131 -1124 9366 -1088
rect 9131 -1144 9299 -1124
rect 7842 -1178 8313 -1159
rect 7789 -1214 8313 -1178
rect 7789 -1219 7957 -1214
rect 6804 -1238 7957 -1219
rect 6804 -1248 6996 -1238
rect 26 -1272 6996 -1248
rect 7030 -1272 7086 -1238
rect 7120 -1272 7176 -1238
rect 7210 -1272 7266 -1238
rect 7300 -1272 7356 -1238
rect 7390 -1272 7446 -1238
rect 7480 -1272 7536 -1238
rect 7570 -1272 7626 -1238
rect 7660 -1272 7716 -1238
rect 7750 -1248 7957 -1238
rect 7991 -1248 8112 -1214
rect 8146 -1219 8313 -1214
rect 9131 -1178 9150 -1144
rect 9184 -1158 9299 -1144
rect 9333 -1158 9366 -1124
rect 9184 -1178 9366 -1158
rect 9131 -1214 9366 -1178
rect 9131 -1219 9299 -1214
rect 8146 -1238 9299 -1219
rect 8146 -1248 8338 -1238
rect 7750 -1272 8338 -1248
rect 8372 -1272 8428 -1238
rect 8462 -1272 8518 -1238
rect 8552 -1272 8608 -1238
rect 8642 -1272 8698 -1238
rect 8732 -1272 8788 -1238
rect 8822 -1272 8878 -1238
rect 8912 -1272 8968 -1238
rect 9002 -1272 9058 -1238
rect 9092 -1248 9299 -1238
rect 9333 -1248 9366 -1214
rect 9092 -1272 9366 -1248
rect 26 -1304 9366 -1272
rect 26 -1338 6770 -1304
rect 6804 -1338 7957 -1304
rect 7991 -1338 8112 -1304
rect 8146 -1338 9299 -1304
rect 9333 -1338 9366 -1304
rect 26 -1388 9366 -1338
rect 26 -1422 6866 -1388
rect 6900 -1422 6956 -1388
rect 6990 -1422 7046 -1388
rect 7080 -1422 7136 -1388
rect 7170 -1422 7226 -1388
rect 7260 -1422 7316 -1388
rect 7350 -1422 7406 -1388
rect 7440 -1422 7496 -1388
rect 7530 -1422 7586 -1388
rect 7620 -1422 7676 -1388
rect 7710 -1422 7766 -1388
rect 7800 -1422 7856 -1388
rect 7890 -1422 8208 -1388
rect 8242 -1422 8298 -1388
rect 8332 -1422 8388 -1388
rect 8422 -1422 8478 -1388
rect 8512 -1422 8568 -1388
rect 8602 -1422 8658 -1388
rect 8692 -1422 8748 -1388
rect 8782 -1422 8838 -1388
rect 8872 -1422 8928 -1388
rect 8962 -1422 9018 -1388
rect 9052 -1422 9108 -1388
rect 9142 -1422 9198 -1388
rect 9232 -1422 9366 -1388
rect 26 -1454 9366 -1422
<< viali >>
rect 379 3825 965 3838
rect 379 3791 426 3825
rect 426 3791 460 3825
rect 460 3791 516 3825
rect 516 3791 550 3825
rect 550 3791 606 3825
rect 606 3791 640 3825
rect 640 3791 696 3825
rect 696 3791 730 3825
rect 730 3791 786 3825
rect 786 3791 820 3825
rect 820 3791 876 3825
rect 876 3791 910 3825
rect 910 3791 965 3825
rect 379 3678 965 3791
rect 379 3644 410 3678
rect 410 3644 444 3678
rect 444 3644 500 3678
rect 500 3644 534 3678
rect 534 3644 590 3678
rect 590 3644 624 3678
rect 624 3644 680 3678
rect 680 3644 714 3678
rect 714 3644 770 3678
rect 770 3644 804 3678
rect 804 3644 860 3678
rect 860 3644 894 3678
rect 894 3644 950 3678
rect 950 3644 965 3678
rect 379 3639 965 3644
<< metal1 >>
rect 360 3838 982 3850
rect 360 3639 379 3838
rect 965 3639 982 3838
rect 360 3514 982 3639
rect 8417 3514 9029 3517
rect 360 2916 9029 3514
rect 360 2781 982 2916
rect 364 -497 976 2781
rect 3047 2181 3661 2184
rect 7076 2182 7690 2184
rect 1702 1546 3664 2181
rect 5732 2174 7690 2182
rect 4463 2092 4941 2122
rect 4463 1644 4474 2092
rect 4924 1644 4941 2092
rect 5729 2110 7690 2174
rect 5729 1630 5808 2110
rect 6262 1630 7690 2110
rect 5729 1546 7690 1630
rect 1704 1436 2318 1546
rect 3047 1436 3661 1546
rect 5729 1436 6343 1546
rect 7076 1436 7690 1546
rect 1703 930 7690 1436
rect 1704 861 2318 930
rect 3047 861 3661 930
rect 1704 227 3661 861
rect 5729 856 6343 930
rect 7076 856 7690 930
rect 1706 225 3661 227
rect 5729 231 7690 856
rect 5729 221 7686 231
rect 5731 220 7686 221
rect 8417 -497 9029 2916
rect 364 -1116 9029 -497
rect 8417 -1118 9029 -1116
<< via1 >>
rect 4474 1644 4924 2092
rect 5808 1630 6262 2110
rect 4458 289 4929 777
<< metal2 >>
rect -234 2092 5008 2188
rect -234 1644 4474 2092
rect 4924 1644 5008 2092
rect -234 1580 5008 1644
rect 5728 2110 9620 2186
rect 5728 1630 5808 2110
rect 6262 1630 9620 2110
rect 5728 1540 9620 1630
rect 4389 777 9658 840
rect 4389 289 4458 777
rect 4929 289 9658 777
rect 4389 228 9658 289
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 ~/share/pdk/sky130A/libs.ref/sky130_fd_pr/mag
timestamp 1746986264
transform 1 0 0 0 1 -138
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1746986264
transform 1 0 1342 0 1 -138
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1746986264
transform 1 0 2684 0 1 -138
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1746986264
transform 1 0 4026 0 1 -138
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1746986264
transform 1 0 5368 0 1 -138
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1746986264
transform 1 0 0 0 1 -1480
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1746986264
transform 1 0 1342 0 1 -1480
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1746986264
transform 1 0 2684 0 1 -1480
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1746986264
transform 1 0 4026 0 1 -1480
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_9
timestamp 1746986264
transform 1 0 5368 0 1 -1480
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_10
timestamp 1746986264
transform 1 0 5368 0 1 2546
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_11
timestamp 1746986264
transform 1 0 4026 0 1 2546
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_12
timestamp 1746986264
transform 1 0 2684 0 1 2546
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_13
timestamp 1746986264
transform 1 0 1342 0 1 2546
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_14
timestamp 1746986264
transform 1 0 0 0 1 2546
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_15
timestamp 1746986264
transform 1 0 5368 0 1 1204
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_16
timestamp 1746986264
transform 1 0 4026 0 1 1204
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17
timestamp 1746986264
transform 1 0 2684 0 1 1204
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_18
timestamp 1746986264
transform 1 0 1342 0 1 1204
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_19
timestamp 1746986264
transform 1 0 0 0 1 1204
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_20
timestamp 1746986264
transform 1 0 6710 0 1 -1480
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_21
timestamp 1746986264
transform 1 0 6710 0 1 -138
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_22
timestamp 1746986264
transform 1 0 8052 0 1 -138
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23
timestamp 1746986264
transform 1 0 8052 0 1 -1480
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_24
timestamp 1746986264
transform 1 0 8052 0 1 1204
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25
timestamp 1746986264
transform 1 0 8052 0 1 2546
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_26
timestamp 1746986264
transform 1 0 6710 0 1 1204
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_27
timestamp 1746986264
transform 1 0 6710 0 1 2546
box 0 0 1340 1340
<< end >>
